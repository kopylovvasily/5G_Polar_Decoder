package pkg;

  //constants responsible for the main Decoder Module
	parameter int BITWIDTH_LLRS = 7;
	parameter int BITWIDTH_REL_SEQ = 10; 
	parameter int N = 512;
	parameter int NR_PROCESSING_UNITS = 64;
  

endpackage


