//This module is used in order to store all the required files that are needed in order to compute the reliability pattern
//The storage is done in a form of Lookup Tables and basicall

module memory_Frozen (
  input logic [2:0] N_i, 
  input logic [5:0] index_i,
  output logic[511:0] Jn_row_o, //only a particular row from the Interleaved Sequence is choosen according to the index
  output logic [511:0][9:0] Jn_Sequence_o,
  output logic [511:0][9:0] Reliability_Sequence_o
);


  logic [511:0][9:0] jn_512;
  logic [255:0][9:0] jn_256;
  logic [127:0][9:0] jn_128;
  logic [63:0][9:0] jn_64;
  logic [31:0][9:0] jn_32;
  logic [511:0][9:0] Reliability_Sequence_512;
  logic [255:0][9:0] Reliability_Sequence_256;
  logic [127:0][9:0] Reliability_Sequence_128;
  logic [63:0][9:0] Reliability_Sequence_64;
  logic [31:0][9:0] Reliability_Sequence_32;
  logic [511:0] row_table_512_o;
  logic [255:0] row_table_256_o;
  logic [127:0] row_table_128_o;
  logic [63:0] row_table_64_o;
  logic [31:0] row_table_32_o;

  //Jn stands for the interleaved Sequence and it is in accrodance with Matworks Notation

  /*************************************************************************************
                          Jn_512
  *************************************************************************************/    

  assign jn_512[511]=10'b0000000000;
  assign jn_512[510]=10'b0000000001;
  assign jn_512[509]=10'b0000000010;
  assign jn_512[508]=10'b0000000011;
  assign jn_512[507]=10'b0000000100;
  assign jn_512[506]=10'b0000000101;
  assign jn_512[505]=10'b0000000110;
  assign jn_512[504]=10'b0000000111;
  assign jn_512[503]=10'b0000001000;
  assign jn_512[502]=10'b0000001001;
  assign jn_512[501]=10'b0000001010;
  assign jn_512[500]=10'b0000001011;
  assign jn_512[499]=10'b0000001100;
  assign jn_512[498]=10'b0000001101;
  assign jn_512[497]=10'b0000001110;
  assign jn_512[496]=10'b0000001111;
  assign jn_512[495]=10'b0000010000;
  assign jn_512[494]=10'b0000010001;
  assign jn_512[493]=10'b0000010010;
  assign jn_512[492]=10'b0000010011;
  assign jn_512[491]=10'b0000010100;
  assign jn_512[490]=10'b0000010101;
  assign jn_512[489]=10'b0000010110;
  assign jn_512[488]=10'b0000010111;
  assign jn_512[487]=10'b0000011000;
  assign jn_512[486]=10'b0000011001;
  assign jn_512[485]=10'b0000011010;
  assign jn_512[484]=10'b0000011011;
  assign jn_512[483]=10'b0000011100;
  assign jn_512[482]=10'b0000011101;
  assign jn_512[481]=10'b0000011110;
  assign jn_512[480]=10'b0000011111;
  assign jn_512[479]=10'b0000100000;
  assign jn_512[478]=10'b0000100001;
  assign jn_512[477]=10'b0000100010;
  assign jn_512[476]=10'b0000100011;
  assign jn_512[475]=10'b0000100100;
  assign jn_512[474]=10'b0000100101;
  assign jn_512[473]=10'b0000100110;
  assign jn_512[472]=10'b0000100111;
  assign jn_512[471]=10'b0000101000;
  assign jn_512[470]=10'b0000101001;
  assign jn_512[469]=10'b0000101010;
  assign jn_512[468]=10'b0000101011;
  assign jn_512[467]=10'b0000101100;
  assign jn_512[466]=10'b0000101101;
  assign jn_512[465]=10'b0000101110;
  assign jn_512[464]=10'b0000101111;
  assign jn_512[463]=10'b0001000000;
  assign jn_512[462]=10'b0001000001;
  assign jn_512[461]=10'b0001000010;
  assign jn_512[460]=10'b0001000011;
  assign jn_512[459]=10'b0001000100;
  assign jn_512[458]=10'b0001000101;
  assign jn_512[457]=10'b0001000110;
  assign jn_512[456]=10'b0001000111;
  assign jn_512[455]=10'b0001001000;
  assign jn_512[454]=10'b0001001001;
  assign jn_512[453]=10'b0001001010;
  assign jn_512[452]=10'b0001001011;
  assign jn_512[451]=10'b0001001100;
  assign jn_512[450]=10'b0001001101;
  assign jn_512[449]=10'b0001001110;
  assign jn_512[448]=10'b0001001111;
  assign jn_512[447]=10'b0000110000;
  assign jn_512[446]=10'b0000110001;
  assign jn_512[445]=10'b0000110010;
  assign jn_512[444]=10'b0000110011;
  assign jn_512[443]=10'b0000110100;
  assign jn_512[442]=10'b0000110101;
  assign jn_512[441]=10'b0000110110;
  assign jn_512[440]=10'b0000110111;
  assign jn_512[439]=10'b0000111000;
  assign jn_512[438]=10'b0000111001;
  assign jn_512[437]=10'b0000111010;
  assign jn_512[436]=10'b0000111011;
  assign jn_512[435]=10'b0000111100;
  assign jn_512[434]=10'b0000111101;
  assign jn_512[433]=10'b0000111110;
  assign jn_512[432]=10'b0000111111;
  assign jn_512[431]=10'b0001010000;
  assign jn_512[430]=10'b0001010001;
  assign jn_512[429]=10'b0001010010;
  assign jn_512[428]=10'b0001010011;
  assign jn_512[427]=10'b0001010100;
  assign jn_512[426]=10'b0001010101;
  assign jn_512[425]=10'b0001010110;
  assign jn_512[424]=10'b0001010111;
  assign jn_512[423]=10'b0001011000;
  assign jn_512[422]=10'b0001011001;
  assign jn_512[421]=10'b0001011010;
  assign jn_512[420]=10'b0001011011;
  assign jn_512[419]=10'b0001011100;
  assign jn_512[418]=10'b0001011101;
  assign jn_512[417]=10'b0001011110;
  assign jn_512[416]=10'b0001011111;
  assign jn_512[415]=10'b0001100000;
  assign jn_512[414]=10'b0001100001;
  assign jn_512[413]=10'b0001100010;
  assign jn_512[412]=10'b0001100011;
  assign jn_512[411]=10'b0001100100;
  assign jn_512[410]=10'b0001100101;
  assign jn_512[409]=10'b0001100110;
  assign jn_512[408]=10'b0001100111;
  assign jn_512[407]=10'b0001101000;
  assign jn_512[406]=10'b0001101001;
  assign jn_512[405]=10'b0001101010;
  assign jn_512[404]=10'b0001101011;
  assign jn_512[403]=10'b0001101100;
  assign jn_512[402]=10'b0001101101;
  assign jn_512[401]=10'b0001101110;
  assign jn_512[400]=10'b0001101111;
  assign jn_512[399]=10'b0001110000;
  assign jn_512[398]=10'b0001110001;
  assign jn_512[397]=10'b0001110010;
  assign jn_512[396]=10'b0001110011;
  assign jn_512[395]=10'b0001110100;
  assign jn_512[394]=10'b0001110101;
  assign jn_512[393]=10'b0001110110;
  assign jn_512[392]=10'b0001110111;
  assign jn_512[391]=10'b0001111000;
  assign jn_512[390]=10'b0001111001;
  assign jn_512[389]=10'b0001111010;
  assign jn_512[388]=10'b0001111011;
  assign jn_512[387]=10'b0001111100;
  assign jn_512[386]=10'b0001111101;
  assign jn_512[385]=10'b0001111110;
  assign jn_512[384]=10'b0001111111;
  assign jn_512[383]=10'b0010000000;
  assign jn_512[382]=10'b0010000001;
  assign jn_512[381]=10'b0010000010;
  assign jn_512[380]=10'b0010000011;
  assign jn_512[379]=10'b0010000100;
  assign jn_512[378]=10'b0010000101;
  assign jn_512[377]=10'b0010000110;
  assign jn_512[376]=10'b0010000111;
  assign jn_512[375]=10'b0010001000;
  assign jn_512[374]=10'b0010001001;
  assign jn_512[373]=10'b0010001010;
  assign jn_512[372]=10'b0010001011;
  assign jn_512[371]=10'b0010001100;
  assign jn_512[370]=10'b0010001101;
  assign jn_512[369]=10'b0010001110;
  assign jn_512[368]=10'b0010001111;
  assign jn_512[367]=10'b0100000000;
  assign jn_512[366]=10'b0100000001;
  assign jn_512[365]=10'b0100000010;
  assign jn_512[364]=10'b0100000011;
  assign jn_512[363]=10'b0100000100;
  assign jn_512[362]=10'b0100000101;
  assign jn_512[361]=10'b0100000110;
  assign jn_512[360]=10'b0100000111;
  assign jn_512[359]=10'b0100001000;
  assign jn_512[358]=10'b0100001001;
  assign jn_512[357]=10'b0100001010;
  assign jn_512[356]=10'b0100001011;
  assign jn_512[355]=10'b0100001100;
  assign jn_512[354]=10'b0100001101;
  assign jn_512[353]=10'b0100001110;
  assign jn_512[352]=10'b0100001111;
  assign jn_512[351]=10'b0010010000;
  assign jn_512[350]=10'b0010010001;
  assign jn_512[349]=10'b0010010010;
  assign jn_512[348]=10'b0010010011;
  assign jn_512[347]=10'b0010010100;
  assign jn_512[346]=10'b0010010101;
  assign jn_512[345]=10'b0010010110;
  assign jn_512[344]=10'b0010010111;
  assign jn_512[343]=10'b0010011000;
  assign jn_512[342]=10'b0010011001;
  assign jn_512[341]=10'b0010011010;
  assign jn_512[340]=10'b0010011011;
  assign jn_512[339]=10'b0010011100;
  assign jn_512[338]=10'b0010011101;
  assign jn_512[337]=10'b0010011110;
  assign jn_512[336]=10'b0010011111;
  assign jn_512[335]=10'b0100010000;
  assign jn_512[334]=10'b0100010001;
  assign jn_512[333]=10'b0100010010;
  assign jn_512[332]=10'b0100010011;
  assign jn_512[331]=10'b0100010100;
  assign jn_512[330]=10'b0100010101;
  assign jn_512[329]=10'b0100010110;
  assign jn_512[328]=10'b0100010111;
  assign jn_512[327]=10'b0100011000;
  assign jn_512[326]=10'b0100011001;
  assign jn_512[325]=10'b0100011010;
  assign jn_512[324]=10'b0100011011;
  assign jn_512[323]=10'b0100011100;
  assign jn_512[322]=10'b0100011101;
  assign jn_512[321]=10'b0100011110;
  assign jn_512[320]=10'b0100011111;
  assign jn_512[319]=10'b0010100000;
  assign jn_512[318]=10'b0010100001;
  assign jn_512[317]=10'b0010100010;
  assign jn_512[316]=10'b0010100011;
  assign jn_512[315]=10'b0010100100;
  assign jn_512[314]=10'b0010100101;
  assign jn_512[313]=10'b0010100110;
  assign jn_512[312]=10'b0010100111;
  assign jn_512[311]=10'b0010101000;
  assign jn_512[310]=10'b0010101001;
  assign jn_512[309]=10'b0010101010;
  assign jn_512[308]=10'b0010101011;
  assign jn_512[307]=10'b0010101100;
  assign jn_512[306]=10'b0010101101;
  assign jn_512[305]=10'b0010101110;
  assign jn_512[304]=10'b0010101111;
  assign jn_512[303]=10'b0100100000;
  assign jn_512[302]=10'b0100100001;
  assign jn_512[301]=10'b0100100010;
  assign jn_512[300]=10'b0100100011;
  assign jn_512[299]=10'b0100100100;
  assign jn_512[298]=10'b0100100101;
  assign jn_512[297]=10'b0100100110;
  assign jn_512[296]=10'b0100100111;
  assign jn_512[295]=10'b0100101000;
  assign jn_512[294]=10'b0100101001;
  assign jn_512[293]=10'b0100101010;
  assign jn_512[292]=10'b0100101011;
  assign jn_512[291]=10'b0100101100;
  assign jn_512[290]=10'b0100101101;
  assign jn_512[289]=10'b0100101110;
  assign jn_512[288]=10'b0100101111;
  assign jn_512[287]=10'b0010110000;
  assign jn_512[286]=10'b0010110001;
  assign jn_512[285]=10'b0010110010;
  assign jn_512[284]=10'b0010110011;
  assign jn_512[283]=10'b0010110100;
  assign jn_512[282]=10'b0010110101;
  assign jn_512[281]=10'b0010110110;
  assign jn_512[280]=10'b0010110111;
  assign jn_512[279]=10'b0010111000;
  assign jn_512[278]=10'b0010111001;
  assign jn_512[277]=10'b0010111010;
  assign jn_512[276]=10'b0010111011;
  assign jn_512[275]=10'b0010111100;
  assign jn_512[274]=10'b0010111101;
  assign jn_512[273]=10'b0010111110;
  assign jn_512[272]=10'b0010111111;
  assign jn_512[271]=10'b0100110000;
  assign jn_512[270]=10'b0100110001;
  assign jn_512[269]=10'b0100110010;
  assign jn_512[268]=10'b0100110011;
  assign jn_512[267]=10'b0100110100;
  assign jn_512[266]=10'b0100110101;
  assign jn_512[265]=10'b0100110110;
  assign jn_512[264]=10'b0100110111;
  assign jn_512[263]=10'b0100111000;
  assign jn_512[262]=10'b0100111001;
  assign jn_512[261]=10'b0100111010;
  assign jn_512[260]=10'b0100111011;
  assign jn_512[259]=10'b0100111100;
  assign jn_512[258]=10'b0100111101;
  assign jn_512[257]=10'b0100111110;
  assign jn_512[256]=10'b0100111111;
  assign jn_512[255]=10'b0011000000;
  assign jn_512[254]=10'b0011000001;
  assign jn_512[253]=10'b0011000010;
  assign jn_512[252]=10'b0011000011;
  assign jn_512[251]=10'b0011000100;
  assign jn_512[250]=10'b0011000101;
  assign jn_512[249]=10'b0011000110;
  assign jn_512[248]=10'b0011000111;
  assign jn_512[247]=10'b0011001000;
  assign jn_512[246]=10'b0011001001;
  assign jn_512[245]=10'b0011001010;
  assign jn_512[244]=10'b0011001011;
  assign jn_512[243]=10'b0011001100;
  assign jn_512[242]=10'b0011001101;
  assign jn_512[241]=10'b0011001110;
  assign jn_512[240]=10'b0011001111;
  assign jn_512[239]=10'b0101000000;
  assign jn_512[238]=10'b0101000001;
  assign jn_512[237]=10'b0101000010;
  assign jn_512[236]=10'b0101000011;
  assign jn_512[235]=10'b0101000100;
  assign jn_512[234]=10'b0101000101;
  assign jn_512[233]=10'b0101000110;
  assign jn_512[232]=10'b0101000111;
  assign jn_512[231]=10'b0101001000;
  assign jn_512[230]=10'b0101001001;
  assign jn_512[229]=10'b0101001010;
  assign jn_512[228]=10'b0101001011;
  assign jn_512[227]=10'b0101001100;
  assign jn_512[226]=10'b0101001101;
  assign jn_512[225]=10'b0101001110;
  assign jn_512[224]=10'b0101001111;
  assign jn_512[223]=10'b0011010000;
  assign jn_512[222]=10'b0011010001;
  assign jn_512[221]=10'b0011010010;
  assign jn_512[220]=10'b0011010011;
  assign jn_512[219]=10'b0011010100;
  assign jn_512[218]=10'b0011010101;
  assign jn_512[217]=10'b0011010110;
  assign jn_512[216]=10'b0011010111;
  assign jn_512[215]=10'b0011011000;
  assign jn_512[214]=10'b0011011001;
  assign jn_512[213]=10'b0011011010;
  assign jn_512[212]=10'b0011011011;
  assign jn_512[211]=10'b0011011100;
  assign jn_512[210]=10'b0011011101;
  assign jn_512[209]=10'b0011011110;
  assign jn_512[208]=10'b0011011111;
  assign jn_512[207]=10'b0101010000;
  assign jn_512[206]=10'b0101010001;
  assign jn_512[205]=10'b0101010010;
  assign jn_512[204]=10'b0101010011;
  assign jn_512[203]=10'b0101010100;
  assign jn_512[202]=10'b0101010101;
  assign jn_512[201]=10'b0101010110;
  assign jn_512[200]=10'b0101010111;
  assign jn_512[199]=10'b0101011000;
  assign jn_512[198]=10'b0101011001;
  assign jn_512[197]=10'b0101011010;
  assign jn_512[196]=10'b0101011011;
  assign jn_512[195]=10'b0101011100;
  assign jn_512[194]=10'b0101011101;
  assign jn_512[193]=10'b0101011110;
  assign jn_512[192]=10'b0101011111;
  assign jn_512[191]=10'b0011100000;
  assign jn_512[190]=10'b0011100001;
  assign jn_512[189]=10'b0011100010;
  assign jn_512[188]=10'b0011100011;
  assign jn_512[187]=10'b0011100100;
  assign jn_512[186]=10'b0011100101;
  assign jn_512[185]=10'b0011100110;
  assign jn_512[184]=10'b0011100111;
  assign jn_512[183]=10'b0011101000;
  assign jn_512[182]=10'b0011101001;
  assign jn_512[181]=10'b0011101010;
  assign jn_512[180]=10'b0011101011;
  assign jn_512[179]=10'b0011101100;
  assign jn_512[178]=10'b0011101101;
  assign jn_512[177]=10'b0011101110;
  assign jn_512[176]=10'b0011101111;
  assign jn_512[175]=10'b0101100000;
  assign jn_512[174]=10'b0101100001;
  assign jn_512[173]=10'b0101100010;
  assign jn_512[172]=10'b0101100011;
  assign jn_512[171]=10'b0101100100;
  assign jn_512[170]=10'b0101100101;
  assign jn_512[169]=10'b0101100110;
  assign jn_512[168]=10'b0101100111;
  assign jn_512[167]=10'b0101101000;
  assign jn_512[166]=10'b0101101001;
  assign jn_512[165]=10'b0101101010;
  assign jn_512[164]=10'b0101101011;
  assign jn_512[163]=10'b0101101100;
  assign jn_512[162]=10'b0101101101;
  assign jn_512[161]=10'b0101101110;
  assign jn_512[160]=10'b0101101111;
  assign jn_512[159]=10'b0011110000;
  assign jn_512[158]=10'b0011110001;
  assign jn_512[157]=10'b0011110010;
  assign jn_512[156]=10'b0011110011;
  assign jn_512[155]=10'b0011110100;
  assign jn_512[154]=10'b0011110101;
  assign jn_512[153]=10'b0011110110;
  assign jn_512[152]=10'b0011110111;
  assign jn_512[151]=10'b0011111000;
  assign jn_512[150]=10'b0011111001;
  assign jn_512[149]=10'b0011111010;
  assign jn_512[148]=10'b0011111011;
  assign jn_512[147]=10'b0011111100;
  assign jn_512[146]=10'b0011111101;
  assign jn_512[145]=10'b0011111110;
  assign jn_512[144]=10'b0011111111;
  assign jn_512[143]=10'b0101110000;
  assign jn_512[142]=10'b0101110001;
  assign jn_512[141]=10'b0101110010;
  assign jn_512[140]=10'b0101110011;
  assign jn_512[139]=10'b0101110100;
  assign jn_512[138]=10'b0101110101;
  assign jn_512[137]=10'b0101110110;
  assign jn_512[136]=10'b0101110111;
  assign jn_512[135]=10'b0101111000;
  assign jn_512[134]=10'b0101111001;
  assign jn_512[133]=10'b0101111010;
  assign jn_512[132]=10'b0101111011;
  assign jn_512[131]=10'b0101111100;
  assign jn_512[130]=10'b0101111101;
  assign jn_512[129]=10'b0101111110;
  assign jn_512[128]=10'b0101111111;
  assign jn_512[127]=10'b0110000000;
  assign jn_512[126]=10'b0110000001;
  assign jn_512[125]=10'b0110000010;
  assign jn_512[124]=10'b0110000011;
  assign jn_512[123]=10'b0110000100;
  assign jn_512[122]=10'b0110000101;
  assign jn_512[121]=10'b0110000110;
  assign jn_512[120]=10'b0110000111;
  assign jn_512[119]=10'b0110001000;
  assign jn_512[118]=10'b0110001001;
  assign jn_512[117]=10'b0110001010;
  assign jn_512[116]=10'b0110001011;
  assign jn_512[115]=10'b0110001100;
  assign jn_512[114]=10'b0110001101;
  assign jn_512[113]=10'b0110001110;
  assign jn_512[112]=10'b0110001111;
  assign jn_512[111]=10'b0110010000;
  assign jn_512[110]=10'b0110010001;
  assign jn_512[109]=10'b0110010010;
  assign jn_512[108]=10'b0110010011;
  assign jn_512[107]=10'b0110010100;
  assign jn_512[106]=10'b0110010101;
  assign jn_512[105]=10'b0110010110;
  assign jn_512[104]=10'b0110010111;
  assign jn_512[103]=10'b0110011000;
  assign jn_512[102]=10'b0110011001;
  assign jn_512[101]=10'b0110011010;
  assign jn_512[100]=10'b0110011011;
  assign jn_512[99]=10'b0110011100;
  assign jn_512[98]=10'b0110011101;
  assign jn_512[97]=10'b0110011110;
  assign jn_512[96]=10'b0110011111;
  assign jn_512[95]=10'b0110100000;
  assign jn_512[94]=10'b0110100001;
  assign jn_512[93]=10'b0110100010;
  assign jn_512[92]=10'b0110100011;
  assign jn_512[91]=10'b0110100100;
  assign jn_512[90]=10'b0110100101;
  assign jn_512[89]=10'b0110100110;
  assign jn_512[88]=10'b0110100111;
  assign jn_512[87]=10'b0110101000;
  assign jn_512[86]=10'b0110101001;
  assign jn_512[85]=10'b0110101010;
  assign jn_512[84]=10'b0110101011;
  assign jn_512[83]=10'b0110101100;
  assign jn_512[82]=10'b0110101101;
  assign jn_512[81]=10'b0110101110;
  assign jn_512[80]=10'b0110101111;
  assign jn_512[79]=10'b0111000000;
  assign jn_512[78]=10'b0111000001;
  assign jn_512[77]=10'b0111000010;
  assign jn_512[76]=10'b0111000011;
  assign jn_512[75]=10'b0111000100;
  assign jn_512[74]=10'b0111000101;
  assign jn_512[73]=10'b0111000110;
  assign jn_512[72]=10'b0111000111;
  assign jn_512[71]=10'b0111001000;
  assign jn_512[70]=10'b0111001001;
  assign jn_512[69]=10'b0111001010;
  assign jn_512[68]=10'b0111001011;
  assign jn_512[67]=10'b0111001100;
  assign jn_512[66]=10'b0111001101;
  assign jn_512[65]=10'b0111001110;
  assign jn_512[64]=10'b0111001111;
  assign jn_512[63]=10'b0110110000;
  assign jn_512[62]=10'b0110110001;
  assign jn_512[61]=10'b0110110010;
  assign jn_512[60]=10'b0110110011;
  assign jn_512[59]=10'b0110110100;
  assign jn_512[58]=10'b0110110101;
  assign jn_512[57]=10'b0110110110;
  assign jn_512[56]=10'b0110110111;
  assign jn_512[55]=10'b0110111000;
  assign jn_512[54]=10'b0110111001;
  assign jn_512[53]=10'b0110111010;
  assign jn_512[52]=10'b0110111011;
  assign jn_512[51]=10'b0110111100;
  assign jn_512[50]=10'b0110111101;
  assign jn_512[49]=10'b0110111110;
  assign jn_512[48]=10'b0110111111;
  assign jn_512[47]=10'b0111010000;
  assign jn_512[46]=10'b0111010001;
  assign jn_512[45]=10'b0111010010;
  assign jn_512[44]=10'b0111010011;
  assign jn_512[43]=10'b0111010100;
  assign jn_512[42]=10'b0111010101;
  assign jn_512[41]=10'b0111010110;
  assign jn_512[40]=10'b0111010111;
  assign jn_512[39]=10'b0111011000;
  assign jn_512[38]=10'b0111011001;
  assign jn_512[37]=10'b0111011010;
  assign jn_512[36]=10'b0111011011;
  assign jn_512[35]=10'b0111011100;
  assign jn_512[34]=10'b0111011101;
  assign jn_512[33]=10'b0111011110;
  assign jn_512[32]=10'b0111011111;
  assign jn_512[31]=10'b0111100000;
  assign jn_512[30]=10'b0111100001;
  assign jn_512[29]=10'b0111100010;
  assign jn_512[28]=10'b0111100011;
  assign jn_512[27]=10'b0111100100;
  assign jn_512[26]=10'b0111100101;
  assign jn_512[25]=10'b0111100110;
  assign jn_512[24]=10'b0111100111;
  assign jn_512[23]=10'b0111101000;
  assign jn_512[22]=10'b0111101001;
  assign jn_512[21]=10'b0111101010;
  assign jn_512[20]=10'b0111101011;
  assign jn_512[19]=10'b0111101100;
  assign jn_512[18]=10'b0111101101;
  assign jn_512[17]=10'b0111101110;
  assign jn_512[16]=10'b0111101111;
  assign jn_512[15]=10'b0111110000;
  assign jn_512[14]=10'b0111110001;
  assign jn_512[13]=10'b0111110010;
  assign jn_512[12]=10'b0111110011;
  assign jn_512[11]=10'b0111110100;
  assign jn_512[10]=10'b0111110101;
  assign jn_512[9]=10'b0111110110;
  assign jn_512[8]=10'b0111110111;
  assign jn_512[7]=10'b0111111000;
  assign jn_512[6]=10'b0111111001;
  assign jn_512[5]=10'b0111111010;
  assign jn_512[4]=10'b0111111011;
  assign jn_512[3]=10'b0111111100;
  assign jn_512[2]=10'b0111111101;
  assign jn_512[1]=10'b0111111110;
  assign jn_512[0]=10'b0111111111;


  /*************************************************************************************
                          Jn_32
  *************************************************************************************/    

  assign jn_32[31]=10'b0000000000;
  assign jn_32[30]=10'b0000000001;
  assign jn_32[29]=10'b0000000010;
  assign jn_32[28]=10'b0000000100;
  assign jn_32[27]=10'b0000000011;
  assign jn_32[26]=10'b0000000101;
  assign jn_32[25]=10'b0000000110;
  assign jn_32[24]=10'b0000000111;
  assign jn_32[23]=10'b0000001000;
  assign jn_32[22]=10'b0000010000;
  assign jn_32[21]=10'b0000001001;
  assign jn_32[20]=10'b0000010001;
  assign jn_32[19]=10'b0000001010;
  assign jn_32[18]=10'b0000010010;
  assign jn_32[17]=10'b0000001011;
  assign jn_32[16]=10'b0000010011;
  assign jn_32[15]=10'b0000001100;
  assign jn_32[14]=10'b0000010100;
  assign jn_32[13]=10'b0000001101;
  assign jn_32[12]=10'b0000010101;
  assign jn_32[11]=10'b0000001110;
  assign jn_32[10]=10'b0000010110;
  assign jn_32[9]=10'b0000001111;
  assign jn_32[8]=10'b0000010111;
  assign jn_32[7]=10'b0000011000;
  assign jn_32[6]=10'b0000011001;
  assign jn_32[5]=10'b0000011010;
  assign jn_32[4]=10'b0000011100;
  assign jn_32[3]=10'b0000011011;
  assign jn_32[2]=10'b0000011101;
  assign jn_32[1]=10'b0000011110;
  assign jn_32[0]=10'b0000011111;

  /*************************************************************************************
                          Jn_64
  *************************************************************************************/    
  assign jn_64[63]=10'b0000000000;
  assign jn_64[62]=10'b0000000001;
  assign jn_64[61]=10'b0000000010;
  assign jn_64[60]=10'b0000000011;
  assign jn_64[59]=10'b0000000100;
  assign jn_64[58]=10'b0000000101;
  assign jn_64[57]=10'b0000001000;
  assign jn_64[56]=10'b0000001001;
  assign jn_64[55]=10'b0000000110;
  assign jn_64[54]=10'b0000000111;
  assign jn_64[53]=10'b0000001010;
  assign jn_64[52]=10'b0000001011;
  assign jn_64[51]=10'b0000001100;
  assign jn_64[50]=10'b0000001101;
  assign jn_64[49]=10'b0000001110;
  assign jn_64[48]=10'b0000001111;
  assign jn_64[47]=10'b0000010000;
  assign jn_64[46]=10'b0000010001;
  assign jn_64[45]=10'b0000100000;
  assign jn_64[44]=10'b0000100001;
  assign jn_64[43]=10'b0000010010;
  assign jn_64[42]=10'b0000010011;
  assign jn_64[41]=10'b0000100010;
  assign jn_64[40]=10'b0000100011;
  assign jn_64[39]=10'b0000010100;
  assign jn_64[38]=10'b0000010101;
  assign jn_64[37]=10'b0000100100;
  assign jn_64[36]=10'b0000100101;
  assign jn_64[35]=10'b0000010110;
  assign jn_64[34]=10'b0000010111;
  assign jn_64[33]=10'b0000100110;
  assign jn_64[32]=10'b0000100111;
  assign jn_64[31]=10'b0000011000;
  assign jn_64[30]=10'b0000011001;
  assign jn_64[29]=10'b0000101000;
  assign jn_64[28]=10'b0000101001;
  assign jn_64[27]=10'b0000011010;
  assign jn_64[26]=10'b0000011011;
  assign jn_64[25]=10'b0000101010;
  assign jn_64[24]=10'b0000101011;
  assign jn_64[23]=10'b0000011100;
  assign jn_64[22]=10'b0000011101;
  assign jn_64[21]=10'b0000101100;
  assign jn_64[20]=10'b0000101101;
  assign jn_64[19]=10'b0000011110;
  assign jn_64[18]=10'b0000011111;
  assign jn_64[17]=10'b0000101110;
  assign jn_64[16]=10'b0000101111;
  assign jn_64[15]=10'b0000110000;
  assign jn_64[14]=10'b0000110001;
  assign jn_64[13]=10'b0000110010;
  assign jn_64[12]=10'b0000110011;
  assign jn_64[11]=10'b0000110100;
  assign jn_64[10]=10'b0000110101;
  assign jn_64[9]=10'b0000111000;
  assign jn_64[8]=10'b0000111001;
  assign jn_64[7]=10'b0000110110;
  assign jn_64[6]=10'b0000110111;
  assign jn_64[5]=10'b0000111010;
  assign jn_64[4]=10'b0000111011;
  assign jn_64[3]=10'b0000111100;
  assign jn_64[2]=10'b0000111101;
  assign jn_64[1]=10'b0000111110;
  assign jn_64[0]=10'b0000111111;

  /*************************************************************************************
                          Jn_128
  *************************************************************************************/    
  assign jn_128[127]=10'b0000000000;
  assign jn_128[126]=10'b0000000001;
  assign jn_128[125]=10'b0000000010;
  assign jn_128[124]=10'b0000000011;
  assign jn_128[123]=10'b0000000100;
  assign jn_128[122]=10'b0000000101;
  assign jn_128[121]=10'b0000000110;
  assign jn_128[120]=10'b0000000111;
  assign jn_128[119]=10'b0000001000;
  assign jn_128[118]=10'b0000001001;
  assign jn_128[117]=10'b0000001010;
  assign jn_128[116]=10'b0000001011;
  assign jn_128[115]=10'b0000010000;
  assign jn_128[114]=10'b0000010001;
  assign jn_128[113]=10'b0000010010;
  assign jn_128[112]=10'b0000010011;
  assign jn_128[111]=10'b0000001100;
  assign jn_128[110]=10'b0000001101;
  assign jn_128[109]=10'b0000001110;
  assign jn_128[108]=10'b0000001111;
  assign jn_128[107]=10'b0000010100;
  assign jn_128[106]=10'b0000010101;
  assign jn_128[105]=10'b0000010110;
  assign jn_128[104]=10'b0000010111;
  assign jn_128[103]=10'b0000011000;
  assign jn_128[102]=10'b0000011001;
  assign jn_128[101]=10'b0000011010;
  assign jn_128[100]=10'b0000011011;
  assign jn_128[99]=10'b0000011100;
  assign jn_128[98]=10'b0000011101;
  assign jn_128[97]=10'b0000011110;
  assign jn_128[96]=10'b0000011111;
  assign jn_128[95]=10'b0000100000;
  assign jn_128[94]=10'b0000100001;
  assign jn_128[93]=10'b0000100010;
  assign jn_128[92]=10'b0000100011;
  assign jn_128[91]=10'b0001000000;
  assign jn_128[90]=10'b0001000001;
  assign jn_128[89]=10'b0001000010;
  assign jn_128[88]=10'b0001000011;
  assign jn_128[87]=10'b0000100100;
  assign jn_128[86]=10'b0000100101;
  assign jn_128[85]=10'b0000100110;
  assign jn_128[84]=10'b0000100111;
  assign jn_128[83]=10'b0001000100;
  assign jn_128[82]=10'b0001000101;
  assign jn_128[81]=10'b0001000110;
  assign jn_128[80]=10'b0001000111;
  assign jn_128[79]=10'b0000101000;
  assign jn_128[78]=10'b0000101001;
  assign jn_128[77]=10'b0000101010;
  assign jn_128[76]=10'b0000101011;
  assign jn_128[75]=10'b0001001000;
  assign jn_128[74]=10'b0001001001;
  assign jn_128[73]=10'b0001001010;
  assign jn_128[72]=10'b0001001011;
  assign jn_128[71]=10'b0000101100;
  assign jn_128[70]=10'b0000101101;
  assign jn_128[69]=10'b0000101110;
  assign jn_128[68]=10'b0000101111;
  assign jn_128[67]=10'b0001001100;
  assign jn_128[66]=10'b0001001101;
  assign jn_128[65]=10'b0001001110;
  assign jn_128[64]=10'b0001001111;
  assign jn_128[63]=10'b0000110000;
  assign jn_128[62]=10'b0000110001;
  assign jn_128[61]=10'b0000110010;
  assign jn_128[60]=10'b0000110011;
  assign jn_128[59]=10'b0001010000;
  assign jn_128[58]=10'b0001010001;
  assign jn_128[57]=10'b0001010010;
  assign jn_128[56]=10'b0001010011;
  assign jn_128[55]=10'b0000110100;
  assign jn_128[54]=10'b0000110101;
  assign jn_128[53]=10'b0000110110;
  assign jn_128[52]=10'b0000110111;
  assign jn_128[51]=10'b0001010100;
  assign jn_128[50]=10'b0001010101;
  assign jn_128[49]=10'b0001010110;
  assign jn_128[48]=10'b0001010111;
  assign jn_128[47]=10'b0000111000;
  assign jn_128[46]=10'b0000111001;
  assign jn_128[45]=10'b0000111010;
  assign jn_128[44]=10'b0000111011;
  assign jn_128[43]=10'b0001011000;
  assign jn_128[42]=10'b0001011001;
  assign jn_128[41]=10'b0001011010;
  assign jn_128[40]=10'b0001011011;
  assign jn_128[39]=10'b0000111100;
  assign jn_128[38]=10'b0000111101;
  assign jn_128[37]=10'b0000111110;
  assign jn_128[36]=10'b0000111111;
  assign jn_128[35]=10'b0001011100;
  assign jn_128[34]=10'b0001011101;
  assign jn_128[33]=10'b0001011110;
  assign jn_128[32]=10'b0001011111;
  assign jn_128[31]=10'b0001100000;
  assign jn_128[30]=10'b0001100001;
  assign jn_128[29]=10'b0001100010;
  assign jn_128[28]=10'b0001100011;
  assign jn_128[27]=10'b0001100100;
  assign jn_128[26]=10'b0001100101;
  assign jn_128[25]=10'b0001100110;
  assign jn_128[24]=10'b0001100111;
  assign jn_128[23]=10'b0001101000;
  assign jn_128[22]=10'b0001101001;
  assign jn_128[21]=10'b0001101010;
  assign jn_128[20]=10'b0001101011;
  assign jn_128[19]=10'b0001110000;
  assign jn_128[18]=10'b0001110001;
  assign jn_128[17]=10'b0001110010;
  assign jn_128[16]=10'b0001110011;
  assign jn_128[15]=10'b0001101100;
  assign jn_128[14]=10'b0001101101;
  assign jn_128[13]=10'b0001101110;
  assign jn_128[12]=10'b0001101111;
  assign jn_128[11]=10'b0001110100;
  assign jn_128[10]=10'b0001110101;
  assign jn_128[9]=10'b0001110110;
  assign jn_128[8]=10'b0001110111;
  assign jn_128[7]=10'b0001111000;
  assign jn_128[6]=10'b0001111001;
  assign jn_128[5]=10'b0001111010;
  assign jn_128[4]=10'b0001111011;
  assign jn_128[3]=10'b0001111100;
  assign jn_128[2]=10'b0001111101;
  assign jn_128[1]=10'b0001111110;
  assign jn_128[0]=10'b0001111111;


  /*************************************************************************************
                          Jn_256
  *************************************************************************************/    
  assign jn_256[255]=10'b0000000000;
  assign jn_256[254]=10'b0000000001;
  assign jn_256[253]=10'b0000000010;
  assign jn_256[252]=10'b0000000011;
  assign jn_256[251]=10'b0000000100;
  assign jn_256[250]=10'b0000000101;
  assign jn_256[249]=10'b0000000110;
  assign jn_256[248]=10'b0000000111;
  assign jn_256[247]=10'b0000001000;
  assign jn_256[246]=10'b0000001001;
  assign jn_256[245]=10'b0000001010;
  assign jn_256[244]=10'b0000001011;
  assign jn_256[243]=10'b0000001100;
  assign jn_256[242]=10'b0000001101;
  assign jn_256[241]=10'b0000001110;
  assign jn_256[240]=10'b0000001111;
  assign jn_256[239]=10'b0000010000;
  assign jn_256[238]=10'b0000010001;
  assign jn_256[237]=10'b0000010010;
  assign jn_256[236]=10'b0000010011;
  assign jn_256[235]=10'b0000010100;
  assign jn_256[234]=10'b0000010101;
  assign jn_256[233]=10'b0000010110;
  assign jn_256[232]=10'b0000010111;
  assign jn_256[231]=10'b0000100000;
  assign jn_256[230]=10'b0000100001;
  assign jn_256[229]=10'b0000100010;
  assign jn_256[228]=10'b0000100011;
  assign jn_256[227]=10'b0000100100;
  assign jn_256[226]=10'b0000100101;
  assign jn_256[225]=10'b0000100110;
  assign jn_256[224]=10'b0000100111;
  assign jn_256[223]=10'b0000011000;
  assign jn_256[222]=10'b0000011001;
  assign jn_256[221]=10'b0000011010;
  assign jn_256[220]=10'b0000011011;
  assign jn_256[219]=10'b0000011100;
  assign jn_256[218]=10'b0000011101;
  assign jn_256[217]=10'b0000011110;
  assign jn_256[216]=10'b0000011111;
  assign jn_256[215]=10'b0000101000;
  assign jn_256[214]=10'b0000101001;
  assign jn_256[213]=10'b0000101010;
  assign jn_256[212]=10'b0000101011;
  assign jn_256[211]=10'b0000101100;
  assign jn_256[210]=10'b0000101101;
  assign jn_256[209]=10'b0000101110;
  assign jn_256[208]=10'b0000101111;
  assign jn_256[207]=10'b0000110000;
  assign jn_256[206]=10'b0000110001;
  assign jn_256[205]=10'b0000110010;
  assign jn_256[204]=10'b0000110011;
  assign jn_256[203]=10'b0000110100;
  assign jn_256[202]=10'b0000110101;
  assign jn_256[201]=10'b0000110110;
  assign jn_256[200]=10'b0000110111;
  assign jn_256[199]=10'b0000111000;
  assign jn_256[198]=10'b0000111001;
  assign jn_256[197]=10'b0000111010;
  assign jn_256[196]=10'b0000111011;
  assign jn_256[195]=10'b0000111100;
  assign jn_256[194]=10'b0000111101;
  assign jn_256[193]=10'b0000111110;
  assign jn_256[192]=10'b0000111111;
  assign jn_256[191]=10'b0001000000;
  assign jn_256[190]=10'b0001000001;
  assign jn_256[189]=10'b0001000010;
  assign jn_256[188]=10'b0001000011;
  assign jn_256[187]=10'b0001000100;
  assign jn_256[186]=10'b0001000101;
  assign jn_256[185]=10'b0001000110;
  assign jn_256[184]=10'b0001000111;
  assign jn_256[183]=10'b0010000000;
  assign jn_256[182]=10'b0010000001;
  assign jn_256[181]=10'b0010000010;
  assign jn_256[180]=10'b0010000011;
  assign jn_256[179]=10'b0010000100;
  assign jn_256[178]=10'b0010000101;
  assign jn_256[177]=10'b0010000110;
  assign jn_256[176]=10'b0010000111;
  assign jn_256[175]=10'b0001001000;
  assign jn_256[174]=10'b0001001001;
  assign jn_256[173]=10'b0001001010;
  assign jn_256[172]=10'b0001001011;
  assign jn_256[171]=10'b0001001100;
  assign jn_256[170]=10'b0001001101;
  assign jn_256[169]=10'b0001001110;
  assign jn_256[168]=10'b0001001111;
  assign jn_256[167]=10'b0010001000;
  assign jn_256[166]=10'b0010001001;
  assign jn_256[165]=10'b0010001010;
  assign jn_256[164]=10'b0010001011;
  assign jn_256[163]=10'b0010001100;
  assign jn_256[162]=10'b0010001101;
  assign jn_256[161]=10'b0010001110;
  assign jn_256[160]=10'b0010001111;
  assign jn_256[159]=10'b0001010000;
  assign jn_256[158]=10'b0001010001;
  assign jn_256[157]=10'b0001010010;
  assign jn_256[156]=10'b0001010011;
  assign jn_256[155]=10'b0001010100;
  assign jn_256[154]=10'b0001010101;
  assign jn_256[153]=10'b0001010110;
  assign jn_256[152]=10'b0001010111;
  assign jn_256[151]=10'b0010010000;
  assign jn_256[150]=10'b0010010001;
  assign jn_256[149]=10'b0010010010;
  assign jn_256[148]=10'b0010010011;
  assign jn_256[147]=10'b0010010100;
  assign jn_256[146]=10'b0010010101;
  assign jn_256[145]=10'b0010010110;
  assign jn_256[144]=10'b0010010111;
  assign jn_256[143]=10'b0001011000;
  assign jn_256[142]=10'b0001011001;
  assign jn_256[141]=10'b0001011010;
  assign jn_256[140]=10'b0001011011;
  assign jn_256[139]=10'b0001011100;
  assign jn_256[138]=10'b0001011101;
  assign jn_256[137]=10'b0001011110;
  assign jn_256[136]=10'b0001011111;
  assign jn_256[135]=10'b0010011000;
  assign jn_256[134]=10'b0010011001;
  assign jn_256[133]=10'b0010011010;
  assign jn_256[132]=10'b0010011011;
  assign jn_256[131]=10'b0010011100;
  assign jn_256[130]=10'b0010011101;
  assign jn_256[129]=10'b0010011110;
  assign jn_256[128]=10'b0010011111;
  assign jn_256[127]=10'b0001100000;
  assign jn_256[126]=10'b0001100001;
  assign jn_256[125]=10'b0001100010;
  assign jn_256[124]=10'b0001100011;
  assign jn_256[123]=10'b0001100100;
  assign jn_256[122]=10'b0001100101;
  assign jn_256[121]=10'b0001100110;
  assign jn_256[120]=10'b0001100111;
  assign jn_256[119]=10'b0010100000;
  assign jn_256[118]=10'b0010100001;
  assign jn_256[117]=10'b0010100010;
  assign jn_256[116]=10'b0010100011;
  assign jn_256[115]=10'b0010100100;
  assign jn_256[114]=10'b0010100101;
  assign jn_256[113]=10'b0010100110;
  assign jn_256[112]=10'b0010100111;
  assign jn_256[111]=10'b0001101000;
  assign jn_256[110]=10'b0001101001;
  assign jn_256[109]=10'b0001101010;
  assign jn_256[108]=10'b0001101011;
  assign jn_256[107]=10'b0001101100;
  assign jn_256[106]=10'b0001101101;
  assign jn_256[105]=10'b0001101110;
  assign jn_256[104]=10'b0001101111;
  assign jn_256[103]=10'b0010101000;
  assign jn_256[102]=10'b0010101001;
  assign jn_256[101]=10'b0010101010;
  assign jn_256[100]=10'b0010101011;
  assign jn_256[99]=10'b0010101100;
  assign jn_256[98]=10'b0010101101;
  assign jn_256[97]=10'b0010101110;
  assign jn_256[96]=10'b0010101111;
  assign jn_256[95]=10'b0001110000;
  assign jn_256[94]=10'b0001110001;
  assign jn_256[93]=10'b0001110010;
  assign jn_256[92]=10'b0001110011;
  assign jn_256[91]=10'b0001110100;
  assign jn_256[90]=10'b0001110101;
  assign jn_256[89]=10'b0001110110;
  assign jn_256[88]=10'b0001110111;
  assign jn_256[87]=10'b0010110000;
  assign jn_256[86]=10'b0010110001;
  assign jn_256[85]=10'b0010110010;
  assign jn_256[84]=10'b0010110011;
  assign jn_256[83]=10'b0010110100;
  assign jn_256[82]=10'b0010110101;
  assign jn_256[81]=10'b0010110110;
  assign jn_256[80]=10'b0010110111;
  assign jn_256[79]=10'b0001111000;
  assign jn_256[78]=10'b0001111001;
  assign jn_256[77]=10'b0001111010;
  assign jn_256[76]=10'b0001111011;
  assign jn_256[75]=10'b0001111100;
  assign jn_256[74]=10'b0001111101;
  assign jn_256[73]=10'b0001111110;
  assign jn_256[72]=10'b0001111111;
  assign jn_256[71]=10'b0010111000;
  assign jn_256[70]=10'b0010111001;
  assign jn_256[69]=10'b0010111010;
  assign jn_256[68]=10'b0010111011;
  assign jn_256[67]=10'b0010111100;
  assign jn_256[66]=10'b0010111101;
  assign jn_256[65]=10'b0010111110;
  assign jn_256[64]=10'b0010111111;
  assign jn_256[63]=10'b0011000000;
  assign jn_256[62]=10'b0011000001;
  assign jn_256[61]=10'b0011000010;
  assign jn_256[60]=10'b0011000011;
  assign jn_256[59]=10'b0011000100;
  assign jn_256[58]=10'b0011000101;
  assign jn_256[57]=10'b0011000110;
  assign jn_256[56]=10'b0011000111;
  assign jn_256[55]=10'b0011001000;
  assign jn_256[54]=10'b0011001001;
  assign jn_256[53]=10'b0011001010;
  assign jn_256[52]=10'b0011001011;
  assign jn_256[51]=10'b0011001100;
  assign jn_256[50]=10'b0011001101;
  assign jn_256[49]=10'b0011001110;
  assign jn_256[48]=10'b0011001111;
  assign jn_256[47]=10'b0011010000;
  assign jn_256[46]=10'b0011010001;
  assign jn_256[45]=10'b0011010010;
  assign jn_256[44]=10'b0011010011;
  assign jn_256[43]=10'b0011010100;
  assign jn_256[42]=10'b0011010101;
  assign jn_256[41]=10'b0011010110;
  assign jn_256[40]=10'b0011010111;
  assign jn_256[39]=10'b0011100000;
  assign jn_256[38]=10'b0011100001;
  assign jn_256[37]=10'b0011100010;
  assign jn_256[36]=10'b0011100011;
  assign jn_256[35]=10'b0011100100;
  assign jn_256[34]=10'b0011100101;
  assign jn_256[33]=10'b0011100110;
  assign jn_256[32]=10'b0011100111;
  assign jn_256[31]=10'b0011011000;
  assign jn_256[30]=10'b0011011001;
  assign jn_256[29]=10'b0011011010;
  assign jn_256[28]=10'b0011011011;
  assign jn_256[27]=10'b0011011100;
  assign jn_256[26]=10'b0011011101;
  assign jn_256[25]=10'b0011011110;
  assign jn_256[24]=10'b0011011111;
  assign jn_256[23]=10'b0011101000;
  assign jn_256[22]=10'b0011101001;
  assign jn_256[21]=10'b0011101010;
  assign jn_256[20]=10'b0011101011;
  assign jn_256[19]=10'b0011101100;
  assign jn_256[18]=10'b0011101101;
  assign jn_256[17]=10'b0011101110;
  assign jn_256[16]=10'b0011101111;
  assign jn_256[15]=10'b0011110000;
  assign jn_256[14]=10'b0011110001;
  assign jn_256[13]=10'b0011110010;
  assign jn_256[12]=10'b0011110011;
  assign jn_256[11]=10'b0011110100;
  assign jn_256[10]=10'b0011110101;
  assign jn_256[9]=10'b0011110110;
  assign jn_256[8]=10'b0011110111;
  assign jn_256[7]=10'b0011111000;
  assign jn_256[6]=10'b0011111001;
  assign jn_256[5]=10'b0011111010;
  assign jn_256[4]=10'b0011111011;
  assign jn_256[3]=10'b0011111100;
  assign jn_256[2]=10'b0011111101;
  assign jn_256[1]=10'b0011111110;
  assign jn_256[0]=10'b0011111111;



  /*************************************************************************************
                          Reliability_Sequence_512
  *************************************************************************************/    
  assign Reliability_Sequence_512[511]=10'b0000000000;
  assign Reliability_Sequence_512[510]=10'b0000000001;
  assign Reliability_Sequence_512[509]=10'b0000000010;
  assign Reliability_Sequence_512[508]=10'b0000000100;
  assign Reliability_Sequence_512[507]=10'b0000001000;
  assign Reliability_Sequence_512[506]=10'b0000010000;
  assign Reliability_Sequence_512[505]=10'b0000100000;
  assign Reliability_Sequence_512[504]=10'b0000000011;
  assign Reliability_Sequence_512[503]=10'b0000000101;
  assign Reliability_Sequence_512[502]=10'b0001000000;
  assign Reliability_Sequence_512[501]=10'b0000001001;
  assign Reliability_Sequence_512[500]=10'b0000000110;
  assign Reliability_Sequence_512[499]=10'b0000010001;
  assign Reliability_Sequence_512[498]=10'b0000001010;
  assign Reliability_Sequence_512[497]=10'b0000010010;
  assign Reliability_Sequence_512[496]=10'b0010000000;
  assign Reliability_Sequence_512[495]=10'b0000001100;
  assign Reliability_Sequence_512[494]=10'b0000100001;
  assign Reliability_Sequence_512[493]=10'b0001000001;
  assign Reliability_Sequence_512[492]=10'b0000010100;
  assign Reliability_Sequence_512[491]=10'b0100000000;
  assign Reliability_Sequence_512[490]=10'b0000100010;
  assign Reliability_Sequence_512[489]=10'b0000011000;
  assign Reliability_Sequence_512[488]=10'b0000100100;
  assign Reliability_Sequence_512[487]=10'b0000000111;
  assign Reliability_Sequence_512[486]=10'b0010000001;
  assign Reliability_Sequence_512[485]=10'b0001000010;
  assign Reliability_Sequence_512[484]=10'b0000001011;
  assign Reliability_Sequence_512[483]=10'b0000101000;
  assign Reliability_Sequence_512[482]=10'b0001000100;
  assign Reliability_Sequence_512[481]=10'b0010000010;
  assign Reliability_Sequence_512[480]=10'b0000010011;
  assign Reliability_Sequence_512[479]=10'b0000001101;
  assign Reliability_Sequence_512[478]=10'b0000110000;
  assign Reliability_Sequence_512[477]=10'b0000001110;
  assign Reliability_Sequence_512[476]=10'b0001001000;
  assign Reliability_Sequence_512[475]=10'b0100000001;
  assign Reliability_Sequence_512[474]=10'b0000010101;
  assign Reliability_Sequence_512[473]=10'b0010000100;
  assign Reliability_Sequence_512[472]=10'b0000100011;
  assign Reliability_Sequence_512[471]=10'b0100000010;
  assign Reliability_Sequence_512[470]=10'b0000011010;
  assign Reliability_Sequence_512[469]=10'b0001010000;
  assign Reliability_Sequence_512[468]=10'b0000100101;
  assign Reliability_Sequence_512[467]=10'b0000011001;
  assign Reliability_Sequence_512[466]=10'b0000010110;
  assign Reliability_Sequence_512[465]=10'b0010001000;
  assign Reliability_Sequence_512[464]=10'b0100000100;
  assign Reliability_Sequence_512[463]=10'b0100001000;
  assign Reliability_Sequence_512[462]=10'b0000100110;
  assign Reliability_Sequence_512[461]=10'b0001100000;
  assign Reliability_Sequence_512[460]=10'b0001000011;
  assign Reliability_Sequence_512[459]=10'b0000101001;
  assign Reliability_Sequence_512[458]=10'b0010010000;
  assign Reliability_Sequence_512[457]=10'b0000011100;
  assign Reliability_Sequence_512[456]=10'b0001000101;
  assign Reliability_Sequence_512[455]=10'b0000101010;
  assign Reliability_Sequence_512[454]=10'b0000110001;
  assign Reliability_Sequence_512[453]=10'b0001001010;
  assign Reliability_Sequence_512[452]=10'b0100010000;
  assign Reliability_Sequence_512[451]=10'b0010100000;
  assign Reliability_Sequence_512[450]=10'b0100100000;
  assign Reliability_Sequence_512[449]=10'b0011000000;
  assign Reliability_Sequence_512[448]=10'b0001000110;
  assign Reliability_Sequence_512[447]=10'b0000101100;
  assign Reliability_Sequence_512[446]=10'b0010000011;
  assign Reliability_Sequence_512[445]=10'b0001010001;
  assign Reliability_Sequence_512[444]=10'b0000110010;
  assign Reliability_Sequence_512[443]=10'b0001001001;
  assign Reliability_Sequence_512[442]=10'b0000001111;
  assign Reliability_Sequence_512[441]=10'b0101000000;
  assign Reliability_Sequence_512[440]=10'b0010000101;
  assign Reliability_Sequence_512[439]=10'b0000110100;
  assign Reliability_Sequence_512[438]=10'b0000010111;
  assign Reliability_Sequence_512[437]=10'b0010000110;
  assign Reliability_Sequence_512[436]=10'b0110000000;
  assign Reliability_Sequence_512[435]=10'b0001001100;
  assign Reliability_Sequence_512[434]=10'b0010001001;
  assign Reliability_Sequence_512[433]=10'b0001010010;
  assign Reliability_Sequence_512[432]=10'b0000111000;
  assign Reliability_Sequence_512[431]=10'b0000011011;
  assign Reliability_Sequence_512[430]=10'b0001100001;
  assign Reliability_Sequence_512[429]=10'b0000100111;
  assign Reliability_Sequence_512[428]=10'b0100000011;
  assign Reliability_Sequence_512[427]=10'b0001010100;
  assign Reliability_Sequence_512[426]=10'b0010001010;
  assign Reliability_Sequence_512[425]=10'b0010010001;
  assign Reliability_Sequence_512[424]=10'b0100000101;
  assign Reliability_Sequence_512[423]=10'b0000011101;
  assign Reliability_Sequence_512[422]=10'b0000101011;
  assign Reliability_Sequence_512[421]=10'b0001100010;
  assign Reliability_Sequence_512[420]=10'b0001011000;
  assign Reliability_Sequence_512[419]=10'b0010001100;
  assign Reliability_Sequence_512[418]=10'b0000011110;
  assign Reliability_Sequence_512[417]=10'b0010010010;
  assign Reliability_Sequence_512[416]=10'b0001000111;
  assign Reliability_Sequence_512[415]=10'b0100000110;
  assign Reliability_Sequence_512[414]=10'b0100001001;
  assign Reliability_Sequence_512[413]=10'b0010100001;
  assign Reliability_Sequence_512[412]=10'b0000101101;
  assign Reliability_Sequence_512[411]=10'b0001100100;
  assign Reliability_Sequence_512[410]=10'b0000110011;
  assign Reliability_Sequence_512[409]=10'b0010010100;
  assign Reliability_Sequence_512[408]=10'b0000101110;
  assign Reliability_Sequence_512[407]=10'b0001001011;
  assign Reliability_Sequence_512[406]=10'b0100001010;
  assign Reliability_Sequence_512[405]=10'b0100010001;
  assign Reliability_Sequence_512[404]=10'b0001101000;
  assign Reliability_Sequence_512[403]=10'b0010100010;
  assign Reliability_Sequence_512[402]=10'b0000110101;
  assign Reliability_Sequence_512[401]=10'b0011000001;
  assign Reliability_Sequence_512[400]=10'b0010011000;
  assign Reliability_Sequence_512[399]=10'b0001001101;
  assign Reliability_Sequence_512[398]=10'b0010100100;
  assign Reliability_Sequence_512[397]=10'b0100001100;
  assign Reliability_Sequence_512[396]=10'b0100010010;
  assign Reliability_Sequence_512[395]=10'b0000110110;
  assign Reliability_Sequence_512[394]=10'b0001010011;
  assign Reliability_Sequence_512[393]=10'b0000111001;
  assign Reliability_Sequence_512[392]=10'b0001110000;
  assign Reliability_Sequence_512[391]=10'b0010000111;
  assign Reliability_Sequence_512[390]=10'b0001001110;
  assign Reliability_Sequence_512[389]=10'b0100100001;
  assign Reliability_Sequence_512[388]=10'b0011000010;
  assign Reliability_Sequence_512[387]=10'b0001010101;
  assign Reliability_Sequence_512[386]=10'b0100010100;
  assign Reliability_Sequence_512[385]=10'b0000111010;
  assign Reliability_Sequence_512[384]=10'b0010101000;
  assign Reliability_Sequence_512[383]=10'b0010001011;
  assign Reliability_Sequence_512[382]=10'b0001100011;
  assign Reliability_Sequence_512[381]=10'b0001010110;
  assign Reliability_Sequence_512[380]=10'b0000111100;
  assign Reliability_Sequence_512[379]=10'b0100011000;
  assign Reliability_Sequence_512[378]=10'b0001011001;
  assign Reliability_Sequence_512[377]=10'b0100100010;
  assign Reliability_Sequence_512[376]=10'b0011000100;
  assign Reliability_Sequence_512[375]=10'b0010001101;
  assign Reliability_Sequence_512[374]=10'b0001100101;
  assign Reliability_Sequence_512[373]=10'b0010010011;
  assign Reliability_Sequence_512[372]=10'b0010110000;
  assign Reliability_Sequence_512[371]=10'b0010001110;
  assign Reliability_Sequence_512[370]=10'b0101000001;
  assign Reliability_Sequence_512[369]=10'b0000011111;
  assign Reliability_Sequence_512[368]=10'b0011001000;
  assign Reliability_Sequence_512[367]=10'b0001011010;
  assign Reliability_Sequence_512[366]=10'b0100100100;
  assign Reliability_Sequence_512[365]=10'b0101000010;
  assign Reliability_Sequence_512[364]=10'b0100000111;
  assign Reliability_Sequence_512[363]=10'b0010010101;
  assign Reliability_Sequence_512[362]=10'b0001100110;
  assign Reliability_Sequence_512[361]=10'b0001101001;
  assign Reliability_Sequence_512[360]=10'b0100110000;
  assign Reliability_Sequence_512[359]=10'b0100101000;
  assign Reliability_Sequence_512[358]=10'b0010100011;
  assign Reliability_Sequence_512[357]=10'b0001011100;
  assign Reliability_Sequence_512[356]=10'b0000101111;
  assign Reliability_Sequence_512[355]=10'b0100001011;
  assign Reliability_Sequence_512[354]=10'b0110000001;
  assign Reliability_Sequence_512[353]=10'b0101000100;
  assign Reliability_Sequence_512[352]=10'b0011010000;
  assign Reliability_Sequence_512[351]=10'b0110000010;
  assign Reliability_Sequence_512[350]=10'b0010010110;
  assign Reliability_Sequence_512[349]=10'b0010011001;
  assign Reliability_Sequence_512[348]=10'b0010100101;
  assign Reliability_Sequence_512[347]=10'b0001101010;
  assign Reliability_Sequence_512[346]=10'b0000110111;
  assign Reliability_Sequence_512[345]=10'b0101001000;
  assign Reliability_Sequence_512[344]=10'b0001110001;
  assign Reliability_Sequence_512[343]=10'b0010011010;
  assign Reliability_Sequence_512[342]=10'b0001001111;
  assign Reliability_Sequence_512[341]=10'b0100001101;
  assign Reliability_Sequence_512[340]=10'b0001101100;
  assign Reliability_Sequence_512[339]=10'b0011100000;
  assign Reliability_Sequence_512[338]=10'b0010100110;
  assign Reliability_Sequence_512[337]=10'b0011000011;
  assign Reliability_Sequence_512[336]=10'b0100001110;
  assign Reliability_Sequence_512[335]=10'b0100010011;
  assign Reliability_Sequence_512[334]=10'b0100100011;
  assign Reliability_Sequence_512[333]=10'b0000111011;
  assign Reliability_Sequence_512[332]=10'b0010101001;
  assign Reliability_Sequence_512[331]=10'b0001110010;
  assign Reliability_Sequence_512[330]=10'b0100010101;
  assign Reliability_Sequence_512[329]=10'b0010011100;
  assign Reliability_Sequence_512[328]=10'b0001010111;
  assign Reliability_Sequence_512[327]=10'b0011000101;
  assign Reliability_Sequence_512[326]=10'b0001110100;
  assign Reliability_Sequence_512[325]=10'b0010101010;
  assign Reliability_Sequence_512[324]=10'b0000111101;
  assign Reliability_Sequence_512[323]=10'b0100011001;
  assign Reliability_Sequence_512[322]=10'b0100010110;
  assign Reliability_Sequence_512[321]=10'b0010110001;
  assign Reliability_Sequence_512[320]=10'b0100100101;
  assign Reliability_Sequence_512[319]=10'b0110000100;
  assign Reliability_Sequence_512[318]=10'b0001011011;
  assign Reliability_Sequence_512[317]=10'b0011000110;
  assign Reliability_Sequence_512[316]=10'b0010101100;
  assign Reliability_Sequence_512[315]=10'b0001111000;
  assign Reliability_Sequence_512[314]=10'b0011001001;
  assign Reliability_Sequence_512[313]=10'b0101010000;
  assign Reliability_Sequence_512[312]=10'b0000111110;
  assign Reliability_Sequence_512[311]=10'b0100011010;
  assign Reliability_Sequence_512[310]=10'b0010001111;
  assign Reliability_Sequence_512[309]=10'b0001100111;
  assign Reliability_Sequence_512[308]=10'b0010110010;
  assign Reliability_Sequence_512[307]=10'b0100100110;
  assign Reliability_Sequence_512[306]=10'b0001011101;
  assign Reliability_Sequence_512[305]=10'b0011001010;
  assign Reliability_Sequence_512[304]=10'b0101000011;
  assign Reliability_Sequence_512[303]=10'b0110001000;
  assign Reliability_Sequence_512[302]=10'b0100101001;
  assign Reliability_Sequence_512[301]=10'b0001101011;
  assign Reliability_Sequence_512[300]=10'b0010110100;
  assign Reliability_Sequence_512[299]=10'b0010010111;
  assign Reliability_Sequence_512[298]=10'b0011010001;
  assign Reliability_Sequence_512[297]=10'b0100011100;
  assign Reliability_Sequence_512[296]=10'b0001011110;
  assign Reliability_Sequence_512[295]=10'b0011001100;
  assign Reliability_Sequence_512[294]=10'b0100101010;
  assign Reliability_Sequence_512[293]=10'b0110010000;
  assign Reliability_Sequence_512[292]=10'b0101100000;
  assign Reliability_Sequence_512[291]=10'b0101000101;
  assign Reliability_Sequence_512[290]=10'b0010011011;
  assign Reliability_Sequence_512[289]=10'b0011010010;
  assign Reliability_Sequence_512[288]=10'b0100110001;
  assign Reliability_Sequence_512[287]=10'b0100101100;
  assign Reliability_Sequence_512[286]=10'b0001101101;
  assign Reliability_Sequence_512[285]=10'b0010111000;
  assign Reliability_Sequence_512[284]=10'b0001110011;
  assign Reliability_Sequence_512[283]=10'b0010100111;
  assign Reliability_Sequence_512[282]=10'b0011100001;
  assign Reliability_Sequence_512[281]=10'b0101000110;
  assign Reliability_Sequence_512[280]=10'b0100110010;
  assign Reliability_Sequence_512[279]=10'b0010011101;
  assign Reliability_Sequence_512[278]=10'b0101001001;
  assign Reliability_Sequence_512[277]=10'b0001101110;
  assign Reliability_Sequence_512[276]=10'b0001110101;
  assign Reliability_Sequence_512[275]=10'b0011010100;
  assign Reliability_Sequence_512[274]=10'b0010101011;
  assign Reliability_Sequence_512[273]=10'b0101001010;
  assign Reliability_Sequence_512[272]=10'b0011100010;
  assign Reliability_Sequence_512[271]=10'b0110000011;
  assign Reliability_Sequence_512[270]=10'b0100110100;
  assign Reliability_Sequence_512[269]=10'b0011011000;
  assign Reliability_Sequence_512[268]=10'b0110100000;
  assign Reliability_Sequence_512[267]=10'b0100001111;
  assign Reliability_Sequence_512[266]=10'b0100010111;
  assign Reliability_Sequence_512[265]=10'b0010011110;
  assign Reliability_Sequence_512[264]=10'b0101010001;
  assign Reliability_Sequence_512[263]=10'b0001110110;
  assign Reliability_Sequence_512[262]=10'b0101001100;
  assign Reliability_Sequence_512[261]=10'b0110000101;
  assign Reliability_Sequence_512[260]=10'b0010101101;
  assign Reliability_Sequence_512[259]=10'b0001111001;
  assign Reliability_Sequence_512[258]=10'b0011000111;
  assign Reliability_Sequence_512[257]=10'b0010110011;
  assign Reliability_Sequence_512[256]=10'b0011100100;
  assign Reliability_Sequence_512[255]=10'b0101010010;
  assign Reliability_Sequence_512[254]=10'b0100111000;
  assign Reliability_Sequence_512[253]=10'b0110000110;
  assign Reliability_Sequence_512[252]=10'b0010101110;
  assign Reliability_Sequence_512[251]=10'b0110001001;
  assign Reliability_Sequence_512[250]=10'b0100011011;
  assign Reliability_Sequence_512[249]=10'b0001111010;
  assign Reliability_Sequence_512[248]=10'b0111000000;
  assign Reliability_Sequence_512[247]=10'b0101100001;
  assign Reliability_Sequence_512[246]=10'b0011001011;
  assign Reliability_Sequence_512[245]=10'b0000111111;
  assign Reliability_Sequence_512[244]=10'b0101010100;
  assign Reliability_Sequence_512[243]=10'b0110001010;
  assign Reliability_Sequence_512[242]=10'b0010110101;
  assign Reliability_Sequence_512[241]=10'b0100100111;
  assign Reliability_Sequence_512[240]=10'b0100011101;
  assign Reliability_Sequence_512[239]=10'b0011101000;
  assign Reliability_Sequence_512[238]=10'b0001111100;
  assign Reliability_Sequence_512[237]=10'b0011001101;
  assign Reliability_Sequence_512[236]=10'b0010110110;
  assign Reliability_Sequence_512[235]=10'b0100011110;
  assign Reliability_Sequence_512[234]=10'b0100101011;
  assign Reliability_Sequence_512[233]=10'b0101100010;
  assign Reliability_Sequence_512[232]=10'b0011010011;
  assign Reliability_Sequence_512[231]=10'b0110010001;
  assign Reliability_Sequence_512[230]=10'b0010111001;
  assign Reliability_Sequence_512[229]=10'b0110001100;
  assign Reliability_Sequence_512[228]=10'b0101011000;
  assign Reliability_Sequence_512[227]=10'b0011110000;
  assign Reliability_Sequence_512[226]=10'b0011001110;
  assign Reliability_Sequence_512[225]=10'b0001011111;
  assign Reliability_Sequence_512[224]=10'b0101000111;
  assign Reliability_Sequence_512[223]=10'b0110010010;
  assign Reliability_Sequence_512[222]=10'b0101100100;
  assign Reliability_Sequence_512[221]=10'b0100110011;
  assign Reliability_Sequence_512[220]=10'b0100101101;
  assign Reliability_Sequence_512[219]=10'b0110100001;
  assign Reliability_Sequence_512[218]=10'b0011010101;
  assign Reliability_Sequence_512[217]=10'b0010111010;
  assign Reliability_Sequence_512[216]=10'b0110010100;
  assign Reliability_Sequence_512[215]=10'b0011100011;
  assign Reliability_Sequence_512[214]=10'b0110100010;
  assign Reliability_Sequence_512[213]=10'b0100101110;
  assign Reliability_Sequence_512[212]=10'b0101101000;
  assign Reliability_Sequence_512[211]=10'b0001101111;
  assign Reliability_Sequence_512[210]=10'b0101001011;
  assign Reliability_Sequence_512[209]=10'b0011010110;
  assign Reliability_Sequence_512[208]=10'b0100110101;
  assign Reliability_Sequence_512[207]=10'b0010111100;
  assign Reliability_Sequence_512[206]=10'b0111000001;
  assign Reliability_Sequence_512[205]=10'b0011011001;
  assign Reliability_Sequence_512[204]=10'b0110011000;
  assign Reliability_Sequence_512[203]=10'b0011100101;
  assign Reliability_Sequence_512[202]=10'b0010011111;
  assign Reliability_Sequence_512[201]=10'b0110100100;
  assign Reliability_Sequence_512[200]=10'b0100110110;
  assign Reliability_Sequence_512[199]=10'b0101001101;
  assign Reliability_Sequence_512[198]=10'b0001110111;
  assign Reliability_Sequence_512[197]=10'b0101010011;
  assign Reliability_Sequence_512[196]=10'b0011011010;
  assign Reliability_Sequence_512[195]=10'b0101110000;
  assign Reliability_Sequence_512[194]=10'b0011100110;
  assign Reliability_Sequence_512[193]=10'b0110000111;
  assign Reliability_Sequence_512[192]=10'b0100111001;
  assign Reliability_Sequence_512[191]=10'b0111000010;
  assign Reliability_Sequence_512[190]=10'b0101001110;
  assign Reliability_Sequence_512[189]=10'b0011101001;
  assign Reliability_Sequence_512[188]=10'b0010101111;
  assign Reliability_Sequence_512[187]=10'b0001111011;
  assign Reliability_Sequence_512[186]=10'b0101010101;
  assign Reliability_Sequence_512[185]=10'b0011011100;
  assign Reliability_Sequence_512[184]=10'b0100111010;
  assign Reliability_Sequence_512[183]=10'b0110101000;
  assign Reliability_Sequence_512[182]=10'b0110001011;
  assign Reliability_Sequence_512[181]=10'b0101100011;
  assign Reliability_Sequence_512[180]=10'b0100011111;
  assign Reliability_Sequence_512[179]=10'b0010110111;
  assign Reliability_Sequence_512[178]=10'b0011101010;
  assign Reliability_Sequence_512[177]=10'b0001111101;
  assign Reliability_Sequence_512[176]=10'b0101010110;
  assign Reliability_Sequence_512[175]=10'b0100111100;
  assign Reliability_Sequence_512[174]=10'b0011110001;
  assign Reliability_Sequence_512[173]=10'b0101011001;
  assign Reliability_Sequence_512[172]=10'b0111000100;
  assign Reliability_Sequence_512[171]=10'b0110001101;
  assign Reliability_Sequence_512[170]=10'b0110010011;
  assign Reliability_Sequence_512[169]=10'b0011001111;
  assign Reliability_Sequence_512[168]=10'b0110110000;
  assign Reliability_Sequence_512[167]=10'b0101100101;
  assign Reliability_Sequence_512[166]=10'b0010111011;
  assign Reliability_Sequence_512[165]=10'b0011101100;
  assign Reliability_Sequence_512[164]=10'b0001111110;
  assign Reliability_Sequence_512[163]=10'b0011110010;
  assign Reliability_Sequence_512[162]=10'b0110001110;
  assign Reliability_Sequence_512[161]=10'b0101011010;
  assign Reliability_Sequence_512[160]=10'b0111001000;
  assign Reliability_Sequence_512[159]=10'b0101100110;
  assign Reliability_Sequence_512[158]=10'b0110010101;
  assign Reliability_Sequence_512[157]=10'b0100101111;
  assign Reliability_Sequence_512[156]=10'b0011110100;
  assign Reliability_Sequence_512[155]=10'b0010111101;
  assign Reliability_Sequence_512[154]=10'b0101101001;
  assign Reliability_Sequence_512[153]=10'b0011010111;
  assign Reliability_Sequence_512[152]=10'b0101011100;
  assign Reliability_Sequence_512[151]=10'b0110100011;
  assign Reliability_Sequence_512[150]=10'b0110010110;
  assign Reliability_Sequence_512[149]=10'b0111010000;
  assign Reliability_Sequence_512[148]=10'b0101101010;
  assign Reliability_Sequence_512[147]=10'b0110011001;
  assign Reliability_Sequence_512[146]=10'b0011011011;
  assign Reliability_Sequence_512[145]=10'b0100110111;
  assign Reliability_Sequence_512[144]=10'b0110100101;
  assign Reliability_Sequence_512[143]=10'b0110011010;
  assign Reliability_Sequence_512[142]=10'b0011100111;
  assign Reliability_Sequence_512[141]=10'b0011111000;
  assign Reliability_Sequence_512[140]=10'b0101110001;
  assign Reliability_Sequence_512[139]=10'b0010111110;
  assign Reliability_Sequence_512[138]=10'b0101101100;
  assign Reliability_Sequence_512[137]=10'b0101001111;
  assign Reliability_Sequence_512[136]=10'b0111100000;
  assign Reliability_Sequence_512[135]=10'b0100111011;
  assign Reliability_Sequence_512[134]=10'b0011011101;
  assign Reliability_Sequence_512[133]=10'b0101110010;
  assign Reliability_Sequence_512[132]=10'b0110100110;
  assign Reliability_Sequence_512[131]=10'b0110101001;
  assign Reliability_Sequence_512[130]=10'b0111000011;
  assign Reliability_Sequence_512[129]=10'b0011101011;
  assign Reliability_Sequence_512[128]=10'b0110011100;
  assign Reliability_Sequence_512[127]=10'b0101010111;
  assign Reliability_Sequence_512[126]=10'b0101110100;
  assign Reliability_Sequence_512[125]=10'b0100111101;
  assign Reliability_Sequence_512[124]=10'b0011011110;
  assign Reliability_Sequence_512[123]=10'b0110101010;
  assign Reliability_Sequence_512[122]=10'b0111000101;
  assign Reliability_Sequence_512[121]=10'b0011101101;
  assign Reliability_Sequence_512[120]=10'b0110110001;
  assign Reliability_Sequence_512[119]=10'b0101011011;
  assign Reliability_Sequence_512[118]=10'b0011110011;
  assign Reliability_Sequence_512[117]=10'b0111000110;
  assign Reliability_Sequence_512[116]=10'b0100111110;
  assign Reliability_Sequence_512[115]=10'b0101111000;
  assign Reliability_Sequence_512[114]=10'b0110101100;
  assign Reliability_Sequence_512[113]=10'b0011101110;
  assign Reliability_Sequence_512[112]=10'b0101100111;
  assign Reliability_Sequence_512[111]=10'b0111001001;
  assign Reliability_Sequence_512[110]=10'b0110001111;
  assign Reliability_Sequence_512[109]=10'b0110110010;
  assign Reliability_Sequence_512[108]=10'b0101011101;
  assign Reliability_Sequence_512[107]=10'b0011110101;
  assign Reliability_Sequence_512[106]=10'b0111001010;
  assign Reliability_Sequence_512[105]=10'b0101101011;
  assign Reliability_Sequence_512[104]=10'b0001111111;
  assign Reliability_Sequence_512[103]=10'b0010111111;
  assign Reliability_Sequence_512[102]=10'b0110010111;
  assign Reliability_Sequence_512[101]=10'b0110110100;
  assign Reliability_Sequence_512[100]=10'b0111010001;
  assign Reliability_Sequence_512[99]=10'b0011110110;
  assign Reliability_Sequence_512[98]=10'b0101011110;
  assign Reliability_Sequence_512[97]=10'b0111001100;
  assign Reliability_Sequence_512[96]=10'b0011111001;
  assign Reliability_Sequence_512[95]=10'b0110011011;
  assign Reliability_Sequence_512[94]=10'b0101101101;
  assign Reliability_Sequence_512[93]=10'b0110111000;
  assign Reliability_Sequence_512[92]=10'b0101110110;
  assign Reliability_Sequence_512[91]=10'b0110100111;
  assign Reliability_Sequence_512[90]=10'b0111010010;
  assign Reliability_Sequence_512[89]=10'b0011111010;
  assign Reliability_Sequence_512[88]=10'b0101110011;
  assign Reliability_Sequence_512[87]=10'b0111100001;
  assign Reliability_Sequence_512[86]=10'b0110011101;
  assign Reliability_Sequence_512[85]=10'b0101101110;
  assign Reliability_Sequence_512[84]=10'b0111010100;
  assign Reliability_Sequence_512[83]=10'b0110101101;
  assign Reliability_Sequence_512[82]=10'b0011111100;
  assign Reliability_Sequence_512[81]=10'b0101110101;
  assign Reliability_Sequence_512[80]=10'b0111100010;
  assign Reliability_Sequence_512[79]=10'b0110101011;
  assign Reliability_Sequence_512[78]=10'b0110011110;
  assign Reliability_Sequence_512[77]=10'b0011011111;
  assign Reliability_Sequence_512[76]=10'b0111011000;
  assign Reliability_Sequence_512[75]=10'b0111000111;
  assign Reliability_Sequence_512[74]=10'b0101111001;
  assign Reliability_Sequence_512[73]=10'b0110110011;
  assign Reliability_Sequence_512[72]=10'b0100111111;
  assign Reliability_Sequence_512[71]=10'b0111100100;
  assign Reliability_Sequence_512[70]=10'b0110101110;
  assign Reliability_Sequence_512[69]=10'b0111101000;
  assign Reliability_Sequence_512[68]=10'b0011101111;
  assign Reliability_Sequence_512[67]=10'b0101111010;
  assign Reliability_Sequence_512[66]=10'b0111001011;
  assign Reliability_Sequence_512[65]=10'b0110110101;
  assign Reliability_Sequence_512[64]=10'b0101111100;
  assign Reliability_Sequence_512[63]=10'b0111001101;
  assign Reliability_Sequence_512[62]=10'b0111110000;
  assign Reliability_Sequence_512[61]=10'b0101011111;
  assign Reliability_Sequence_512[60]=10'b0111010011;
  assign Reliability_Sequence_512[59]=10'b0110110110;
  assign Reliability_Sequence_512[58]=10'b0011111011;
  assign Reliability_Sequence_512[57]=10'b0111001110;
  assign Reliability_Sequence_512[56]=10'b0110111010;
  assign Reliability_Sequence_512[55]=10'b0110111001;
  assign Reliability_Sequence_512[54]=10'b0111010101;
  assign Reliability_Sequence_512[53]=10'b0011110111;
  assign Reliability_Sequence_512[52]=10'b0101101111;
  assign Reliability_Sequence_512[51]=10'b0011111101;
  assign Reliability_Sequence_512[50]=10'b0101110111;
  assign Reliability_Sequence_512[49]=10'b0110111100;
  assign Reliability_Sequence_512[48]=10'b0111010110;
  assign Reliability_Sequence_512[47]=10'b0111100011;
  assign Reliability_Sequence_512[46]=10'b0110011111;
  assign Reliability_Sequence_512[45]=10'b0111100101;
  assign Reliability_Sequence_512[44]=10'b0111011001;
  assign Reliability_Sequence_512[43]=10'b0111011010;
  assign Reliability_Sequence_512[42]=10'b0011111110;
  assign Reliability_Sequence_512[41]=10'b0101111011;
  assign Reliability_Sequence_512[40]=10'b0110101111;
  assign Reliability_Sequence_512[39]=10'b0111101001;
  assign Reliability_Sequence_512[38]=10'b0111100110;
  assign Reliability_Sequence_512[37]=10'b0111011100;
  assign Reliability_Sequence_512[36]=10'b0110110111;
  assign Reliability_Sequence_512[35]=10'b0111101010;
  assign Reliability_Sequence_512[34]=10'b0111001111;
  assign Reliability_Sequence_512[33]=10'b0101111101;
  assign Reliability_Sequence_512[32]=10'b0111110001;
  assign Reliability_Sequence_512[31]=10'b0111101100;
  assign Reliability_Sequence_512[30]=10'b0110111011;
  assign Reliability_Sequence_512[29]=10'b0101111110;
  assign Reliability_Sequence_512[28]=10'b0111110010;
  assign Reliability_Sequence_512[27]=10'b0110111101;
  assign Reliability_Sequence_512[26]=10'b0111010111;
  assign Reliability_Sequence_512[25]=10'b0111110100;
  assign Reliability_Sequence_512[24]=10'b0110111110;
  assign Reliability_Sequence_512[23]=10'b0111011011;
  assign Reliability_Sequence_512[22]=10'b0111100111;
  assign Reliability_Sequence_512[21]=10'b0111111000;
  assign Reliability_Sequence_512[20]=10'b0011111111;
  assign Reliability_Sequence_512[19]=10'b0111011101;
  assign Reliability_Sequence_512[18]=10'b0111101011;
  assign Reliability_Sequence_512[17]=10'b0111011110;
  assign Reliability_Sequence_512[16]=10'b0101111111;
  assign Reliability_Sequence_512[15]=10'b0111101101;
  assign Reliability_Sequence_512[14]=10'b0111110011;
  assign Reliability_Sequence_512[13]=10'b0111110110;
  assign Reliability_Sequence_512[12]=10'b0111101110;
  assign Reliability_Sequence_512[11]=10'b0111110101;
  assign Reliability_Sequence_512[10]=10'b0110111111;
  assign Reliability_Sequence_512[9]=10'b0111111001;
  assign Reliability_Sequence_512[8]=10'b0111111010;
  assign Reliability_Sequence_512[7]=10'b0111011111;
  assign Reliability_Sequence_512[6]=10'b0111111100;
  assign Reliability_Sequence_512[5]=10'b0111101111;
  assign Reliability_Sequence_512[4]=10'b0111110111;
  assign Reliability_Sequence_512[3]=10'b0111111011;
  assign Reliability_Sequence_512[2]=10'b0111111101;
  assign Reliability_Sequence_512[1]=10'b0111111110;
  assign Reliability_Sequence_512[0]=10'b0111111111; 


  /*************************************************************************************
                          Reliability_Sequence_32
  *************************************************************************************/    

  assign Reliability_Sequence_32[31]=10'b0000000000;
  assign Reliability_Sequence_32[30]=10'b0000000001;
  assign Reliability_Sequence_32[29]=10'b0000000010;
  assign Reliability_Sequence_32[28]=10'b0000000100;
  assign Reliability_Sequence_32[27]=10'b0000001000;
  assign Reliability_Sequence_32[26]=10'b0000010000;
  assign Reliability_Sequence_32[25]=10'b0000000011;
  assign Reliability_Sequence_32[24]=10'b0000000101;
  assign Reliability_Sequence_32[23]=10'b0000001001;
  assign Reliability_Sequence_32[22]=10'b0000000110;
  assign Reliability_Sequence_32[21]=10'b0000010001;
  assign Reliability_Sequence_32[20]=10'b0000001010;
  assign Reliability_Sequence_32[19]=10'b0000010010;
  assign Reliability_Sequence_32[18]=10'b0000001100;
  assign Reliability_Sequence_32[17]=10'b0000010100;
  assign Reliability_Sequence_32[16]=10'b0000011000;
  assign Reliability_Sequence_32[15]=10'b0000000111;
  assign Reliability_Sequence_32[14]=10'b0000001011;
  assign Reliability_Sequence_32[13]=10'b0000010011;
  assign Reliability_Sequence_32[12]=10'b0000001101;
  assign Reliability_Sequence_32[11]=10'b0000001110;
  assign Reliability_Sequence_32[10]=10'b0000010101;
  assign Reliability_Sequence_32[9]=10'b0000011010;
  assign Reliability_Sequence_32[8]=10'b0000011001;
  assign Reliability_Sequence_32[7]=10'b0000010110;
  assign Reliability_Sequence_32[6]=10'b0000011100;
  assign Reliability_Sequence_32[5]=10'b0000001111;
  assign Reliability_Sequence_32[4]=10'b0000010111;
  assign Reliability_Sequence_32[3]=10'b0000011011;
  assign Reliability_Sequence_32[2]=10'b0000011101;
  assign Reliability_Sequence_32[1]=10'b0000011110;
  assign Reliability_Sequence_32[0]=10'b0000011111;

  /*************************************************************************************
                  Reliability_Sequence_64
  *************************************************************************************/    
  assign Reliability_Sequence_64[63]=10'b0000000000;
  assign Reliability_Sequence_64[62]=10'b0000000001;
  assign Reliability_Sequence_64[61]=10'b0000000010;
  assign Reliability_Sequence_64[60]=10'b0000000100;
  assign Reliability_Sequence_64[59]=10'b0000001000;
  assign Reliability_Sequence_64[58]=10'b0000010000;
  assign Reliability_Sequence_64[57]=10'b0000100000;
  assign Reliability_Sequence_64[56]=10'b0000000011;
  assign Reliability_Sequence_64[55]=10'b0000000101;
  assign Reliability_Sequence_64[54]=10'b0000001001;
  assign Reliability_Sequence_64[53]=10'b0000000110;
  assign Reliability_Sequence_64[52]=10'b0000010001;
  assign Reliability_Sequence_64[51]=10'b0000001010;
  assign Reliability_Sequence_64[50]=10'b0000010010;
  assign Reliability_Sequence_64[49]=10'b0000001100;
  assign Reliability_Sequence_64[48]=10'b0000100001;
  assign Reliability_Sequence_64[47]=10'b0000010100;
  assign Reliability_Sequence_64[46]=10'b0000100010;
  assign Reliability_Sequence_64[45]=10'b0000011000;
  assign Reliability_Sequence_64[44]=10'b0000100100;
  assign Reliability_Sequence_64[43]=10'b0000000111;
  assign Reliability_Sequence_64[42]=10'b0000001011;
  assign Reliability_Sequence_64[41]=10'b0000101000;
  assign Reliability_Sequence_64[40]=10'b0000010011;
  assign Reliability_Sequence_64[39]=10'b0000001101;
  assign Reliability_Sequence_64[38]=10'b0000110000;
  assign Reliability_Sequence_64[37]=10'b0000001110;
  assign Reliability_Sequence_64[36]=10'b0000010101;
  assign Reliability_Sequence_64[35]=10'b0000100011;
  assign Reliability_Sequence_64[34]=10'b0000011010;
  assign Reliability_Sequence_64[33]=10'b0000100101;
  assign Reliability_Sequence_64[32]=10'b0000011001;
  assign Reliability_Sequence_64[31]=10'b0000010110;
  assign Reliability_Sequence_64[30]=10'b0000100110;
  assign Reliability_Sequence_64[29]=10'b0000101001;
  assign Reliability_Sequence_64[28]=10'b0000011100;
  assign Reliability_Sequence_64[27]=10'b0000101010;
  assign Reliability_Sequence_64[26]=10'b0000110001;
  assign Reliability_Sequence_64[25]=10'b0000101100;
  assign Reliability_Sequence_64[24]=10'b0000110010;
  assign Reliability_Sequence_64[23]=10'b0000001111;
  assign Reliability_Sequence_64[22]=10'b0000110100;
  assign Reliability_Sequence_64[21]=10'b0000010111;
  assign Reliability_Sequence_64[20]=10'b0000111000;
  assign Reliability_Sequence_64[19]=10'b0000011011;
  assign Reliability_Sequence_64[18]=10'b0000100111;
  assign Reliability_Sequence_64[17]=10'b0000011101;
  assign Reliability_Sequence_64[16]=10'b0000101011;
  assign Reliability_Sequence_64[15]=10'b0000011110;
  assign Reliability_Sequence_64[14]=10'b0000101101;
  assign Reliability_Sequence_64[13]=10'b0000110011;
  assign Reliability_Sequence_64[12]=10'b0000101110;
  assign Reliability_Sequence_64[11]=10'b0000110101;
  assign Reliability_Sequence_64[10]=10'b0000110110;
  assign Reliability_Sequence_64[9]=10'b0000111001;
  assign Reliability_Sequence_64[8]=10'b0000111010;
  assign Reliability_Sequence_64[7]=10'b0000111100;
  assign Reliability_Sequence_64[6]=10'b0000011111;
  assign Reliability_Sequence_64[5]=10'b0000101111;
  assign Reliability_Sequence_64[4]=10'b0000110111;
  assign Reliability_Sequence_64[3]=10'b0000111011;
  assign Reliability_Sequence_64[2]=10'b0000111101;
  assign Reliability_Sequence_64[1]=10'b0000111110;
  assign Reliability_Sequence_64[0]=10'b0000111111;

  /*************************************************************************************
                  Reliability_Sequence_128
  *************************************************************************************/    

  assign Reliability_Sequence_128[127]=10'b0000000000;
  assign Reliability_Sequence_128[126]=10'b0000000001;
  assign Reliability_Sequence_128[125]=10'b0000000010;
  assign Reliability_Sequence_128[124]=10'b0000000100;
  assign Reliability_Sequence_128[123]=10'b0000001000;
  assign Reliability_Sequence_128[122]=10'b0000010000;
  assign Reliability_Sequence_128[121]=10'b0000100000;
  assign Reliability_Sequence_128[120]=10'b0000000011;
  assign Reliability_Sequence_128[119]=10'b0000000101;
  assign Reliability_Sequence_128[118]=10'b0001000000;
  assign Reliability_Sequence_128[117]=10'b0000001001;
  assign Reliability_Sequence_128[116]=10'b0000000110;
  assign Reliability_Sequence_128[115]=10'b0000010001;
  assign Reliability_Sequence_128[114]=10'b0000001010;
  assign Reliability_Sequence_128[113]=10'b0000010010;
  assign Reliability_Sequence_128[112]=10'b0000001100;
  assign Reliability_Sequence_128[111]=10'b0000100001;
  assign Reliability_Sequence_128[110]=10'b0001000001;
  assign Reliability_Sequence_128[109]=10'b0000010100;
  assign Reliability_Sequence_128[108]=10'b0000100010;
  assign Reliability_Sequence_128[107]=10'b0000011000;
  assign Reliability_Sequence_128[106]=10'b0000100100;
  assign Reliability_Sequence_128[105]=10'b0000000111;
  assign Reliability_Sequence_128[104]=10'b0001000010;
  assign Reliability_Sequence_128[103]=10'b0000001011;
  assign Reliability_Sequence_128[102]=10'b0000101000;
  assign Reliability_Sequence_128[101]=10'b0001000100;
  assign Reliability_Sequence_128[100]=10'b0000010011;
  assign Reliability_Sequence_128[99]=10'b0000001101;
  assign Reliability_Sequence_128[98]=10'b0000110000;
  assign Reliability_Sequence_128[97]=10'b0000001110;
  assign Reliability_Sequence_128[96]=10'b0001001000;
  assign Reliability_Sequence_128[95]=10'b0000010101;
  assign Reliability_Sequence_128[94]=10'b0000100011;
  assign Reliability_Sequence_128[93]=10'b0000011010;
  assign Reliability_Sequence_128[92]=10'b0001010000;
  assign Reliability_Sequence_128[91]=10'b0000100101;
  assign Reliability_Sequence_128[90]=10'b0000011001;
  assign Reliability_Sequence_128[89]=10'b0000010110;
  assign Reliability_Sequence_128[88]=10'b0000100110;
  assign Reliability_Sequence_128[87]=10'b0001100000;
  assign Reliability_Sequence_128[86]=10'b0001000011;
  assign Reliability_Sequence_128[85]=10'b0000101001;
  assign Reliability_Sequence_128[84]=10'b0000011100;
  assign Reliability_Sequence_128[83]=10'b0001000101;
  assign Reliability_Sequence_128[82]=10'b0000101010;
  assign Reliability_Sequence_128[81]=10'b0000110001;
  assign Reliability_Sequence_128[80]=10'b0001001010;
  assign Reliability_Sequence_128[79]=10'b0001000110;
  assign Reliability_Sequence_128[78]=10'b0000101100;
  assign Reliability_Sequence_128[77]=10'b0001010001;
  assign Reliability_Sequence_128[76]=10'b0000110010;
  assign Reliability_Sequence_128[75]=10'b0001001001;
  assign Reliability_Sequence_128[74]=10'b0000001111;
  assign Reliability_Sequence_128[73]=10'b0000110100;
  assign Reliability_Sequence_128[72]=10'b0000010111;
  assign Reliability_Sequence_128[71]=10'b0001001100;
  assign Reliability_Sequence_128[70]=10'b0001010010;
  assign Reliability_Sequence_128[69]=10'b0000111000;
  assign Reliability_Sequence_128[68]=10'b0000011011;
  assign Reliability_Sequence_128[67]=10'b0001100001;
  assign Reliability_Sequence_128[66]=10'b0000100111;
  assign Reliability_Sequence_128[65]=10'b0001010100;
  assign Reliability_Sequence_128[64]=10'b0000011101;
  assign Reliability_Sequence_128[63]=10'b0000101011;
  assign Reliability_Sequence_128[62]=10'b0001100010;
  assign Reliability_Sequence_128[61]=10'b0001011000;
  assign Reliability_Sequence_128[60]=10'b0000011110;
  assign Reliability_Sequence_128[59]=10'b0001000111;
  assign Reliability_Sequence_128[58]=10'b0000101101;
  assign Reliability_Sequence_128[57]=10'b0001100100;
  assign Reliability_Sequence_128[56]=10'b0000110011;
  assign Reliability_Sequence_128[55]=10'b0000101110;
  assign Reliability_Sequence_128[54]=10'b0001001011;
  assign Reliability_Sequence_128[53]=10'b0001101000;
  assign Reliability_Sequence_128[52]=10'b0000110101;
  assign Reliability_Sequence_128[51]=10'b0001001101;
  assign Reliability_Sequence_128[50]=10'b0000110110;
  assign Reliability_Sequence_128[49]=10'b0001010011;
  assign Reliability_Sequence_128[48]=10'b0000111001;
  assign Reliability_Sequence_128[47]=10'b0001110000;
  assign Reliability_Sequence_128[46]=10'b0001001110;
  assign Reliability_Sequence_128[45]=10'b0001010101;
  assign Reliability_Sequence_128[44]=10'b0000111010;
  assign Reliability_Sequence_128[43]=10'b0001100011;
  assign Reliability_Sequence_128[42]=10'b0001010110;
  assign Reliability_Sequence_128[41]=10'b0000111100;
  assign Reliability_Sequence_128[40]=10'b0001011001;
  assign Reliability_Sequence_128[39]=10'b0001100101;
  assign Reliability_Sequence_128[38]=10'b0000011111;
  assign Reliability_Sequence_128[37]=10'b0001011010;
  assign Reliability_Sequence_128[36]=10'b0001100110;
  assign Reliability_Sequence_128[35]=10'b0001101001;
  assign Reliability_Sequence_128[34]=10'b0001011100;
  assign Reliability_Sequence_128[33]=10'b0000101111;
  assign Reliability_Sequence_128[32]=10'b0001101010;
  assign Reliability_Sequence_128[31]=10'b0000110111;
  assign Reliability_Sequence_128[30]=10'b0001110001;
  assign Reliability_Sequence_128[29]=10'b0001001111;
  assign Reliability_Sequence_128[28]=10'b0001101100;
  assign Reliability_Sequence_128[27]=10'b0000111011;
  assign Reliability_Sequence_128[26]=10'b0001110010;
  assign Reliability_Sequence_128[25]=10'b0001010111;
  assign Reliability_Sequence_128[24]=10'b0001110100;
  assign Reliability_Sequence_128[23]=10'b0000111101;
  assign Reliability_Sequence_128[22]=10'b0001011011;
  assign Reliability_Sequence_128[21]=10'b0001111000;
  assign Reliability_Sequence_128[20]=10'b0000111110;
  assign Reliability_Sequence_128[19]=10'b0001100111;
  assign Reliability_Sequence_128[18]=10'b0001011101;
  assign Reliability_Sequence_128[17]=10'b0001101011;
  assign Reliability_Sequence_128[16]=10'b0001011110;
  assign Reliability_Sequence_128[15]=10'b0001101101;
  assign Reliability_Sequence_128[14]=10'b0001110011;
  assign Reliability_Sequence_128[13]=10'b0001101110;
  assign Reliability_Sequence_128[12]=10'b0001110101;
  assign Reliability_Sequence_128[11]=10'b0001110110;
  assign Reliability_Sequence_128[10]=10'b0001111001;
  assign Reliability_Sequence_128[9]=10'b0001111010;
  assign Reliability_Sequence_128[8]=10'b0000111111;
  assign Reliability_Sequence_128[7]=10'b0001111100;
  assign Reliability_Sequence_128[6]=10'b0001011111;
  assign Reliability_Sequence_128[5]=10'b0001101111;
  assign Reliability_Sequence_128[4]=10'b0001110111;
  assign Reliability_Sequence_128[3]=10'b0001111011;
  assign Reliability_Sequence_128[2]=10'b0001111101;
  assign Reliability_Sequence_128[1]=10'b0001111110;
  assign Reliability_Sequence_128[0]=10'b0001111111;

  /*************************************************************************************
                  Reliability_Sequence_256
  *************************************************************************************/    

  assign Reliability_Sequence_256[255]=10'b0000000000;
  assign Reliability_Sequence_256[254]=10'b0000000001;
  assign Reliability_Sequence_256[253]=10'b0000000010;
  assign Reliability_Sequence_256[252]=10'b0000000100;
  assign Reliability_Sequence_256[251]=10'b0000001000;
  assign Reliability_Sequence_256[250]=10'b0000010000;
  assign Reliability_Sequence_256[249]=10'b0000100000;
  assign Reliability_Sequence_256[248]=10'b0000000011;
  assign Reliability_Sequence_256[247]=10'b0000000101;
  assign Reliability_Sequence_256[246]=10'b0001000000;
  assign Reliability_Sequence_256[245]=10'b0000001001;
  assign Reliability_Sequence_256[244]=10'b0000000110;
  assign Reliability_Sequence_256[243]=10'b0000010001;
  assign Reliability_Sequence_256[242]=10'b0000001010;
  assign Reliability_Sequence_256[241]=10'b0000010010;
  assign Reliability_Sequence_256[240]=10'b0010000000;
  assign Reliability_Sequence_256[239]=10'b0000001100;
  assign Reliability_Sequence_256[238]=10'b0000100001;
  assign Reliability_Sequence_256[237]=10'b0001000001;
  assign Reliability_Sequence_256[236]=10'b0000010100;
  assign Reliability_Sequence_256[235]=10'b0000100010;
  assign Reliability_Sequence_256[234]=10'b0000011000;
  assign Reliability_Sequence_256[233]=10'b0000100100;
  assign Reliability_Sequence_256[232]=10'b0000000111;
  assign Reliability_Sequence_256[231]=10'b0010000001;
  assign Reliability_Sequence_256[230]=10'b0001000010;
  assign Reliability_Sequence_256[229]=10'b0000001011;
  assign Reliability_Sequence_256[228]=10'b0000101000;
  assign Reliability_Sequence_256[227]=10'b0001000100;
  assign Reliability_Sequence_256[226]=10'b0010000010;
  assign Reliability_Sequence_256[225]=10'b0000010011;
  assign Reliability_Sequence_256[224]=10'b0000001101;
  assign Reliability_Sequence_256[223]=10'b0000110000;
  assign Reliability_Sequence_256[222]=10'b0000001110;
  assign Reliability_Sequence_256[221]=10'b0001001000;
  assign Reliability_Sequence_256[220]=10'b0000010101;
  assign Reliability_Sequence_256[219]=10'b0010000100;
  assign Reliability_Sequence_256[218]=10'b0000100011;
  assign Reliability_Sequence_256[217]=10'b0000011010;
  assign Reliability_Sequence_256[216]=10'b0001010000;
  assign Reliability_Sequence_256[215]=10'b0000100101;
  assign Reliability_Sequence_256[214]=10'b0000011001;
  assign Reliability_Sequence_256[213]=10'b0000010110;
  assign Reliability_Sequence_256[212]=10'b0010001000;
  assign Reliability_Sequence_256[211]=10'b0000100110;
  assign Reliability_Sequence_256[210]=10'b0001100000;
  assign Reliability_Sequence_256[209]=10'b0001000011;
  assign Reliability_Sequence_256[208]=10'b0000101001;
  assign Reliability_Sequence_256[207]=10'b0010010000;
  assign Reliability_Sequence_256[206]=10'b0000011100;
  assign Reliability_Sequence_256[205]=10'b0001000101;
  assign Reliability_Sequence_256[204]=10'b0000101010;
  assign Reliability_Sequence_256[203]=10'b0000110001;
  assign Reliability_Sequence_256[202]=10'b0001001010;
  assign Reliability_Sequence_256[201]=10'b0010100000;
  assign Reliability_Sequence_256[200]=10'b0011000000;
  assign Reliability_Sequence_256[199]=10'b0001000110;
  assign Reliability_Sequence_256[198]=10'b0000101100;
  assign Reliability_Sequence_256[197]=10'b0010000011;
  assign Reliability_Sequence_256[196]=10'b0001010001;
  assign Reliability_Sequence_256[195]=10'b0000110010;
  assign Reliability_Sequence_256[194]=10'b0001001001;
  assign Reliability_Sequence_256[193]=10'b0000001111;
  assign Reliability_Sequence_256[192]=10'b0010000101;
  assign Reliability_Sequence_256[191]=10'b0000110100;
  assign Reliability_Sequence_256[190]=10'b0000010111;
  assign Reliability_Sequence_256[189]=10'b0010000110;
  assign Reliability_Sequence_256[188]=10'b0001001100;
  assign Reliability_Sequence_256[187]=10'b0010001001;
  assign Reliability_Sequence_256[186]=10'b0001010010;
  assign Reliability_Sequence_256[185]=10'b0000111000;
  assign Reliability_Sequence_256[184]=10'b0000011011;
  assign Reliability_Sequence_256[183]=10'b0001100001;
  assign Reliability_Sequence_256[182]=10'b0000100111;
  assign Reliability_Sequence_256[181]=10'b0001010100;
  assign Reliability_Sequence_256[180]=10'b0010001010;
  assign Reliability_Sequence_256[179]=10'b0010010001;
  assign Reliability_Sequence_256[178]=10'b0000011101;
  assign Reliability_Sequence_256[177]=10'b0000101011;
  assign Reliability_Sequence_256[176]=10'b0001100010;
  assign Reliability_Sequence_256[175]=10'b0001011000;
  assign Reliability_Sequence_256[174]=10'b0010001100;
  assign Reliability_Sequence_256[173]=10'b0000011110;
  assign Reliability_Sequence_256[172]=10'b0010010010;
  assign Reliability_Sequence_256[171]=10'b0001000111;
  assign Reliability_Sequence_256[170]=10'b0010100001;
  assign Reliability_Sequence_256[169]=10'b0000101101;
  assign Reliability_Sequence_256[168]=10'b0001100100;
  assign Reliability_Sequence_256[167]=10'b0000110011;
  assign Reliability_Sequence_256[166]=10'b0010010100;
  assign Reliability_Sequence_256[165]=10'b0000101110;
  assign Reliability_Sequence_256[164]=10'b0001001011;
  assign Reliability_Sequence_256[163]=10'b0001101000;
  assign Reliability_Sequence_256[162]=10'b0010100010;
  assign Reliability_Sequence_256[161]=10'b0000110101;
  assign Reliability_Sequence_256[160]=10'b0011000001;
  assign Reliability_Sequence_256[159]=10'b0010011000;
  assign Reliability_Sequence_256[158]=10'b0001001101;
  assign Reliability_Sequence_256[157]=10'b0010100100;
  assign Reliability_Sequence_256[156]=10'b0000110110;
  assign Reliability_Sequence_256[155]=10'b0001010011;
  assign Reliability_Sequence_256[154]=10'b0000111001;
  assign Reliability_Sequence_256[153]=10'b0001110000;
  assign Reliability_Sequence_256[152]=10'b0010000111;
  assign Reliability_Sequence_256[151]=10'b0001001110;
  assign Reliability_Sequence_256[150]=10'b0011000010;
  assign Reliability_Sequence_256[149]=10'b0001010101;
  assign Reliability_Sequence_256[148]=10'b0000111010;
  assign Reliability_Sequence_256[147]=10'b0010101000;
  assign Reliability_Sequence_256[146]=10'b0010001011;
  assign Reliability_Sequence_256[145]=10'b0001100011;
  assign Reliability_Sequence_256[144]=10'b0001010110;
  assign Reliability_Sequence_256[143]=10'b0000111100;
  assign Reliability_Sequence_256[142]=10'b0001011001;
  assign Reliability_Sequence_256[141]=10'b0011000100;
  assign Reliability_Sequence_256[140]=10'b0010001101;
  assign Reliability_Sequence_256[139]=10'b0001100101;
  assign Reliability_Sequence_256[138]=10'b0010010011;
  assign Reliability_Sequence_256[137]=10'b0010110000;
  assign Reliability_Sequence_256[136]=10'b0010001110;
  assign Reliability_Sequence_256[135]=10'b0000011111;
  assign Reliability_Sequence_256[134]=10'b0011001000;
  assign Reliability_Sequence_256[133]=10'b0001011010;
  assign Reliability_Sequence_256[132]=10'b0010010101;
  assign Reliability_Sequence_256[131]=10'b0001100110;
  assign Reliability_Sequence_256[130]=10'b0001101001;
  assign Reliability_Sequence_256[129]=10'b0010100011;
  assign Reliability_Sequence_256[128]=10'b0001011100;
  assign Reliability_Sequence_256[127]=10'b0000101111;
  assign Reliability_Sequence_256[126]=10'b0011010000;
  assign Reliability_Sequence_256[125]=10'b0010010110;
  assign Reliability_Sequence_256[124]=10'b0010011001;
  assign Reliability_Sequence_256[123]=10'b0010100101;
  assign Reliability_Sequence_256[122]=10'b0001101010;
  assign Reliability_Sequence_256[121]=10'b0000110111;
  assign Reliability_Sequence_256[120]=10'b0001110001;
  assign Reliability_Sequence_256[119]=10'b0010011010;
  assign Reliability_Sequence_256[118]=10'b0001001111;
  assign Reliability_Sequence_256[117]=10'b0001101100;
  assign Reliability_Sequence_256[116]=10'b0011100000;
  assign Reliability_Sequence_256[115]=10'b0010100110;
  assign Reliability_Sequence_256[114]=10'b0011000011;
  assign Reliability_Sequence_256[113]=10'b0000111011;
  assign Reliability_Sequence_256[112]=10'b0010101001;
  assign Reliability_Sequence_256[111]=10'b0001110010;
  assign Reliability_Sequence_256[110]=10'b0010011100;
  assign Reliability_Sequence_256[109]=10'b0001010111;
  assign Reliability_Sequence_256[108]=10'b0011000101;
  assign Reliability_Sequence_256[107]=10'b0001110100;
  assign Reliability_Sequence_256[106]=10'b0010101010;
  assign Reliability_Sequence_256[105]=10'b0000111101;
  assign Reliability_Sequence_256[104]=10'b0010110001;
  assign Reliability_Sequence_256[103]=10'b0001011011;
  assign Reliability_Sequence_256[102]=10'b0011000110;
  assign Reliability_Sequence_256[101]=10'b0010101100;
  assign Reliability_Sequence_256[100]=10'b0001111000;
  assign Reliability_Sequence_256[99]=10'b0011001001;
  assign Reliability_Sequence_256[98]=10'b0000111110;
  assign Reliability_Sequence_256[97]=10'b0010001111;
  assign Reliability_Sequence_256[96]=10'b0001100111;
  assign Reliability_Sequence_256[95]=10'b0010110010;
  assign Reliability_Sequence_256[94]=10'b0001011101;
  assign Reliability_Sequence_256[93]=10'b0011001010;
  assign Reliability_Sequence_256[92]=10'b0001101011;
  assign Reliability_Sequence_256[91]=10'b0010110100;
  assign Reliability_Sequence_256[90]=10'b0010010111;
  assign Reliability_Sequence_256[89]=10'b0011010001;
  assign Reliability_Sequence_256[88]=10'b0001011110;
  assign Reliability_Sequence_256[87]=10'b0011001100;
  assign Reliability_Sequence_256[86]=10'b0010011011;
  assign Reliability_Sequence_256[85]=10'b0011010010;
  assign Reliability_Sequence_256[84]=10'b0001101101;
  assign Reliability_Sequence_256[83]=10'b0010111000;
  assign Reliability_Sequence_256[82]=10'b0001110011;
  assign Reliability_Sequence_256[81]=10'b0010100111;
  assign Reliability_Sequence_256[80]=10'b0011100001;
  assign Reliability_Sequence_256[79]=10'b0010011101;
  assign Reliability_Sequence_256[78]=10'b0001101110;
  assign Reliability_Sequence_256[77]=10'b0001110101;
  assign Reliability_Sequence_256[76]=10'b0011010100;
  assign Reliability_Sequence_256[75]=10'b0010101011;
  assign Reliability_Sequence_256[74]=10'b0011100010;
  assign Reliability_Sequence_256[73]=10'b0011011000;
  assign Reliability_Sequence_256[72]=10'b0010011110;
  assign Reliability_Sequence_256[71]=10'b0001110110;
  assign Reliability_Sequence_256[70]=10'b0010101101;
  assign Reliability_Sequence_256[69]=10'b0001111001;
  assign Reliability_Sequence_256[68]=10'b0011000111;
  assign Reliability_Sequence_256[67]=10'b0010110011;
  assign Reliability_Sequence_256[66]=10'b0011100100;
  assign Reliability_Sequence_256[65]=10'b0010101110;
  assign Reliability_Sequence_256[64]=10'b0001111010;
  assign Reliability_Sequence_256[63]=10'b0011001011;
  assign Reliability_Sequence_256[62]=10'b0000111111;
  assign Reliability_Sequence_256[61]=10'b0010110101;
  assign Reliability_Sequence_256[60]=10'b0011101000;
  assign Reliability_Sequence_256[59]=10'b0001111100;
  assign Reliability_Sequence_256[58]=10'b0011001101;
  assign Reliability_Sequence_256[57]=10'b0010110110;
  assign Reliability_Sequence_256[56]=10'b0011010011;
  assign Reliability_Sequence_256[55]=10'b0010111001;
  assign Reliability_Sequence_256[54]=10'b0011110000;
  assign Reliability_Sequence_256[53]=10'b0011001110;
  assign Reliability_Sequence_256[52]=10'b0001011111;
  assign Reliability_Sequence_256[51]=10'b0011010101;
  assign Reliability_Sequence_256[50]=10'b0010111010;
  assign Reliability_Sequence_256[49]=10'b0011100011;
  assign Reliability_Sequence_256[48]=10'b0001101111;
  assign Reliability_Sequence_256[47]=10'b0011010110;
  assign Reliability_Sequence_256[46]=10'b0010111100;
  assign Reliability_Sequence_256[45]=10'b0011011001;
  assign Reliability_Sequence_256[44]=10'b0011100101;
  assign Reliability_Sequence_256[43]=10'b0010011111;
  assign Reliability_Sequence_256[42]=10'b0001110111;
  assign Reliability_Sequence_256[41]=10'b0011011010;
  assign Reliability_Sequence_256[40]=10'b0011100110;
  assign Reliability_Sequence_256[39]=10'b0011101001;
  assign Reliability_Sequence_256[38]=10'b0010101111;
  assign Reliability_Sequence_256[37]=10'b0001111011;
  assign Reliability_Sequence_256[36]=10'b0011011100;
  assign Reliability_Sequence_256[35]=10'b0010110111;
  assign Reliability_Sequence_256[34]=10'b0011101010;
  assign Reliability_Sequence_256[33]=10'b0001111101;
  assign Reliability_Sequence_256[32]=10'b0011110001;
  assign Reliability_Sequence_256[31]=10'b0011001111;
  assign Reliability_Sequence_256[30]=10'b0010111011;
  assign Reliability_Sequence_256[29]=10'b0011101100;
  assign Reliability_Sequence_256[28]=10'b0001111110;
  assign Reliability_Sequence_256[27]=10'b0011110010;
  assign Reliability_Sequence_256[26]=10'b0011110100;
  assign Reliability_Sequence_256[25]=10'b0010111101;
  assign Reliability_Sequence_256[24]=10'b0011010111;
  assign Reliability_Sequence_256[23]=10'b0011011011;
  assign Reliability_Sequence_256[22]=10'b0011100111;
  assign Reliability_Sequence_256[21]=10'b0011111000;
  assign Reliability_Sequence_256[20]=10'b0010111110;
  assign Reliability_Sequence_256[19]=10'b0011011101;
  assign Reliability_Sequence_256[18]=10'b0011101011;
  assign Reliability_Sequence_256[17]=10'b0011011110;
  assign Reliability_Sequence_256[16]=10'b0011101101;
  assign Reliability_Sequence_256[15]=10'b0011110011;
  assign Reliability_Sequence_256[14]=10'b0011101110;
  assign Reliability_Sequence_256[13]=10'b0011110101;
  assign Reliability_Sequence_256[12]=10'b0001111111;
  assign Reliability_Sequence_256[11]=10'b0010111111;
  assign Reliability_Sequence_256[10]=10'b0011110110;
  assign Reliability_Sequence_256[9]=10'b0011111001;
  assign Reliability_Sequence_256[8]=10'b0011111010;
  assign Reliability_Sequence_256[7]=10'b0011111100;
  assign Reliability_Sequence_256[6]=10'b0011011111;
  assign Reliability_Sequence_256[5]=10'b0011101111;
  assign Reliability_Sequence_256[4]=10'b0011111011;
  assign Reliability_Sequence_256[3]=10'b0011110111;
  assign Reliability_Sequence_256[2]=10'b0011111101;
  assign Reliability_Sequence_256[1]=10'b0011111110;
  assign Reliability_Sequence_256[0]=10'b0011111111;



  always_comb begin
    row_table_512_o = '0;
    row_table_256_o = '0;
    row_table_128_o = '0;
    row_table_64_o = '0;
    row_table_32_o = '0;
    for (int i = 0; i < 512; i++) begin
     Reliability_Sequence_o[i] = 10'b1111111111;
    end
    for (int i = 0; i < 512; i++) begin
     Jn_Sequence_o[i] = 10'b1111111111;
    end 
    Jn_row_o = '0;

    if(N_i == 3'b110) begin //512
      case(index_i)

        6'd0: row_table_512_o = '0;
        6'd1: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000100000000101000000100000000000000101000001100100110010010011001001111101101111111;
        6'd2: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000010000000000000001000000000010000000110000001001001001000100010010101000100101100111000011101110001111100111011111111011101111111111111111;
        6'd3: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000001000010000000100001000000000100000001000000000010001000000010000000010100001000000010001110000001101001001001010010000110010001011001001100110011010111001101101101111000011101110011111110111011111111011101111111111111111;
        6'd4: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000010000000000000001000000000100000000000000000000010010000001000000010100100001000000000001010000010001001010000000101001000000010100000001100000000011101000001010100000011101001100000010001110100001101001001001110010001110010101011001101100111011010111001101101101111000011111110011111110111011111111011101111111111111111;
        6'd5: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000010000000000000001000000000100000000000000000000010010000001000000010100100001000000000001010100010001001010000000101001000001010100000001100000001011101000011010101000011101001101100010011110101001101011011001110110001111011101111111101111111011110111011111101111111101111111111111111111111111111111111111111111111111111;
        6'd6: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000001000000000000000000010000000000000001000000000110000000001000000000110010000001000010010100110001000100000101010100011001001110100000101101000001110101000001110010001011101101011011101010011111001111101010011111101001111011011111110111001111011111111111111111111011110111111111101111111111111111111111111111111111111111111111111111111111111;
        6'd7: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000000001000000000000000000010000010000000001000010000110010000001000000100110110001001000011010100110011000100000111011100011001101110100100111101000111110101001101110010101111101101011111101011111111101111101010111111111011111111011111111111001111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd8: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000000100000001000010000000000000000000000000000000000100000000000010000000000010000010100100000000001111000001000001010000000001000000010100110000000111000010010111010000001100100101110110001011001011010100111011000101000111011110111001101110101100111101010111110111001101110010101111111101011111101011111111101111101110111111111011111111011111111111001111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd9: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000000100000001000010000000000000000000000000000000000100000000000010000000000010001010100100001000001111000001000001010000000001000001010100110000100111001010010111011001001110100101111110001011001111110100111011100101100111111110111101111110101111111101110111111111001111110110111111111111011111101111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd10: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000000000011100000001000010000000000000000000000100000000010100100000000110001000000110001010101100001110001111001001000001110010100001010001110110110000110111101010011111011101011110100111111110001011101111111100111011110101101111111110111111111111101111111101110111111111101111110110111111111111011111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd11: row_table_512_o = 512'b00000000000000000000000000000000000000000000000000000100000111100000001000010000000000100000001000100010001010110101000000110101000010110011010101101001110001111111001010001110110101101010111110110110100110111101111011111111101011111100111111110111011101111111110111011111101111111111110111111111111101111111111110111111111101111111110111111111111011111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd12: row_table_512_o = 512'b00000000000000010000100001000010000010101000001110000100000111100100001100110100000101110000101011100010011010110111000010110101100010111011110101111001110011111111001010101111110101101010111110110110110110111101111011111111101011111100111111111111011101111111110111011111101111111111110111111111111101111111111110111111111101111111110111111111111011111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd13: row_table_512_o = 512'b00000000000000010000100001000010000010101000001110100100000111100100001100110100010101110010101011101010011110110111000110110101110010111111110101111111110011111111101110111111110111101110111110111110111110111111111011111111111111111111111111111111111111111111111111011111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd14: row_table_512_o = 512'b00000000000000010000100001000010010010101010001110100100010111100111001110110111010111110011101011101110011111110111111110111111111111111111110111111111111011111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd15: row_table_512_o = 512'b00000010010000010110110101101110010110111011001111111101111111111111101110111111011111110111101111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd16: row_table_512_o = '0;
        6'd17: row_table_512_o =512'b11111101101111101001001010010001101001000100110000000010000000000000010001000000100000001000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd18: row_table_512_o =512'b11111111111111101111011110111101101101010101110001011011101000011000110001001000101000001100010100010001100000001000000001000000000000000000001000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd19: row_table_512_o =512'b11111111111111101111011110111101111101010111110001011011111000011011110011001011101010001101010100010101100001001000111001001010001101000000001010000000001100000000010001000000001000010001000001000001000001000000000100000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd20: row_table_512_o =512'b11111111111111101111011110111101111101010111110001111011111000011011110011001011111010001111010100011101100101001000111101001010011101000100001010000110001100000000110101010000001010010101000001001001001001000010000100000000010100000011000000000000100010000000001000100000010000000000001000000000000010000000000001000000000010000000001000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd21: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111011111000011111110111101111111111011111110111011101110101001010111111001010111101001100101010010110001110000000110101110001001010010101000001001001011001000010000100000000010100000011000000001000100010000000001000100000010000000000001000000000000010000000000001000000000010000000001000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd22: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111100011111110111101111111111111111111111011111111101011011111111001110111111001110101010011110001110000110110111110001101011110101110001001001111001000010101100000100010100001011000000001110100010000000011000100001010010000000001000000000000010000000010001000000000010000001001000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd23: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111111011111110111101111111111111111111111111111111111011111111111101111111111101110101011011110111110000111110111110101111111110111110101011001111011000110101101000100110110001011010000001110100110000001011000100011010011000000001000010000001010000000010001000000000110000001001000000000000100000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd24: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111111011111110111101111111111111111111111111111111111011111111111101111111111101111101011011111111110000111110111110101111111110111111101011001111111000111101101000101111110011011010001001110100110100101011000100111010111000100001000110010001010011000010101000001000110010001101010000000010100000010100000000010000010001000000000100000000100000000000110000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd25: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111110111111111111111111101111101111111110111101111001101111110111111011001001110110111100101011001100111011111000100011100110010001011011000010111000001010110010001101010000010010100000010100000000010000010101000000000100000000100000000000110000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd26: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111110111111111111111111101111111111111110111111111001111111110111111111001101111110111101101011001110111011111010101011100110110001011111010010111110001010111110001101110100010010100100010101100000110000010101100000010110000100100000001000110000100000000000000000000100001000000000010000000000000000000000000000000000000000000000000000000000000;
        6'd27: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111101111111111111110111111111011111111111111111111101101111110111111101011011110111111111110101011101110110101111111010110111110101011111110011111110100010111100101010111100010110010011101100001010110010100100110001001110000100010000000010000000100001000100000010000000010000000000000000000000000000000000000000000000000000;
        6'd28: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111101111111111111110111111111011111111111111111111101101111110111111101011011110111111111110101111101110110101111111010110111111101011111110011111111100010111110101011111100010110011111101110001011110010110110110001101110001101010100110010011000100101000110010010010000111100000001100000001000100000000100010000000000000000;
        6'd29: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111011111111111111111111111111110111101111111011110111111111011111110111111111101110111111101111111101011110111111101110001111110010110110110101101111001101110100110110011001100101000110010010010000111100010001100000001000100000000100010000000000000000;
        6'd30: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111011111111111101111111111111110111111111101111111001111110110110110111011101101010111011010011000111100010001110000011000100000000100010000000000000000;
        6'd31: row_table_512_o =512'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111110111111011111111010111111011111111111111010111110011011001101101100110110000010010000000;
    
      endcase 

    Reliability_Sequence_o = Reliability_Sequence_512;
    Jn_Sequence_o = jn_512;
    Jn_row_o = row_table_512_o;

    end else if(N_i == 3'b101)begin //256

      case(index_i)
        6'd0: row_table_256_o = '0;  
        6'd1: row_table_256_o = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000001000000001000101001010100101100101011111110011111111111;
        6'd2: row_table_256_o = 256'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000001000000001000000100000001000000000101000001000001001000001000101010000100010110000101001001010101101010101100111001010110101101111011111110011111111111;
        6'd3: row_table_256_o = 256'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000001001000000001000100100000001000001000101001001100101011000101010101010110100110110101111011011111111101110111101111011111111111111111111111111111111111111;
        6'd4: row_table_256_o = 256'b0000000000000000000000000000000000000000000001000000001100000000000000001000000100000101000011010010001001001010001010100100111001001101001111011001110101111001101110101011111101111110111111111011111111101111111101111111111111111111111111111111111111111111;
        6'd5: row_table_256_o = 256'b0000000000000000000000000000000000000001000001001000001100010000000001001010100110010101010011011010101001101011011011100111111101111101101111011111110111111001111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111;
        6'd6: row_table_256_o = 256'b0000000001000001001000001100110000101001000101101010011110110101001111001011100111011101010111011110101111101111011111110111111101111101111111011111110111111011111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111;
        6'd7: row_table_256_o = 256'b0000000001000001001001001101110010101011010101111111111111111101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        6'd8: row_table_256_o = '0;
        6'd9: row_table_256_o = 256'b1111111110111110110110110010001101010100101010000000000000000010010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd10: row_table_256_o = 256'b1111111110111110110111110011001111010110111010010101100001001010110000110100011000100010101000100001010000010000100000001000000010000010000000100000001000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;
        6'd11: row_table_256_o =256'b1111111111111111111111111111111111111110111110110111110011101111111110110101011001101010101100100101010110010100100100011000000010000010010000100000001000000110000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;
        6'd12: row_table_256_o =256'b1111111111111111111111111111111111111111111110111111110011111111111111110111111011111010111100101101110110110101110101011011000110110010110000100110001010000110010001010100000010000001000000000100000000010000000010000000000000000000000000000000000000000000;
        6'd13: row_table_256_o =256'b1111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111101111110110111111110111011011111110111110111010110110011010100111010101010101001011001001010000100100000000010001000010000100000000000000000000000000000000000000;
        6'd14: row_table_256_o =256'b1111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111101111111110111111110111111011111110111111111010111110111110110111110111010101111011101001111010110110101010010101010011000110101001010010000100000001100000000000;
        6'd15: row_table_256_o =256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110111110111111110111010110101011010011010100000001100000000000;
      endcase 

    Reliability_Sequence_o[255:0] = Reliability_Sequence_256;
    Jn_Sequence_o[255:0] = jn_256;
    Jn_row_o[255:0] = row_table_256_o;

    end else if(N_i == 3'b100) begin //128
      case(index_i)

        6'd0: row_table_128_o = '0;
        6'd1: row_table_128_o = 128'b00000000000000000000000000000000000000001000000000000000000010000100001000100000100010001001100101010101001010101111111010111111;
        6'd2: row_table_128_o = 128'b00000000000000000000000000000100000100001000001000110010011010100110001100110111101111111011110111011111111111111111111111111111;
        6'd3: row_table_128_o = 128'b00000010010000001101010101100101010110011110111111111010111011101110111111111111111111111011111111111111111111111111111111111111;
        6'd4: row_table_128_o = '0;
        6'd5: row_table_128_o = 128'b11111101101111110010101010011010101001100001000000000101000100010001000000000000000000000100000000000000000000000000000000000000;
        6'd6: row_table_128_o = 128'b11111111111111111111111111111011111011110111110111001101100101011001110011001000010000000100001000100000000000000000000000000000;
        6'd7: row_table_128_o = 128'b11111111111111111111111111111111111111110111111111111111111101111011110111011111011101110110011010101010110101010000000101000000;      

      endcase 

    Reliability_Sequence_o[127:0] = Reliability_Sequence_128;
    Jn_Sequence_o[127:0] = jn_128;
    Jn_row_o[127:0] = row_table_128_o;

    end else if(N_i == 3'b011) begin //64
      case(index_i)
        6'd0: row_table_64_o = '0;
        6'd1: row_table_64_o = 64'b0000000000000000001000100100010100111111010110111111111111111111;
        6'd2: row_table_64_o = '0;
        6'd3: row_table_64_o = 64'b1111111111111111110111011011101011000000101001000000000000000000;
      endcase 

    Reliability_Sequence_o[63:0] = Reliability_Sequence_64;
    Jn_Sequence_o[63:0] = jn_64;
    Jn_row_o[63:0] = row_table_64_o;

    end else if(N_i == 3'b010) begin //32
      case(index_i)
        6'd0: row_table_32_o = '0;
        6'd1: row_table_32_o = '0;
      endcase 
    Reliability_Sequence_o[31:0] = Reliability_Sequence_32;
    Jn_Sequence_o[31:0] = jn_32;
    Jn_row_o[31:0] = row_table_32_o;
    end
  end
endmodule 